BZh91AY&SY�h�� �_�Px����������`��R�  A�����I!h#M4S��i����L�� jz *!A��@    `�1 �&	�!��L�����Q��   4�  mU�     @  $Ђ	6����O�1�124`&h~�B74@�'`�OAZ�<�a�i6� & ���?�/��HX$x�9'�s���<�z#������q��/�333.���������������� �!�?����Im/]zt������O,�ԦL���8p_T�P�< q2s..U񤡳`̭�yN��lKU�Y���y'����=��m���ؽE�Ъbe�t�n:�+,��A&�8���U�J��'���@���r�6���y��]��/k�K"F��q)(��]�$,I�Y�1�oϾ��##+��4Qۮ�z8E
Zz�-����0�b����!��t��J�״��+ ���g��)[�����a-�2$�&m*m�h@���!ЛL"%d�x��< �@*�D9Nd�� $��I��!÷���� ���ӅS�o��Wm%S����Իl��1�SG��+$���H�b(e����@�q�0ZX�Sj^e�F��ʕ.0��T�KLC P�Y��1��&�юûNq�ݕ���D�l��c���u,�(����B�XtC��U	I��xnkp�~5�\u�y�lϏm����%�޶��V�GH'�j�nXyn�d[�g-p�W)Vaq�Pmn�����U#���Z��j� �<�0`�i8�.���A	n0��J��MM2L�3`�\�A�@ͽJ�L6b1HWʍF�k����wMڭ�Řp�V�9I;ܮ8}�q�iN��zi�WE�^�mCc��u�,�W�qM8�Eȉ��M�)<kv��Z��t6늕�R4at��Ö^J�1����QW����~:��:=*�&�ɠ^������a�7��Ī�"Q$(R$AH�&�ޘ�5��,a$QF&���4���ZF�rܫK���%Kk$�(��M��vZ���h�Uy�Tk=<��$�6bʗ:����z'�Q)�'��Y�h���>Q��i�F�h�	�1>7~�m*Q'���?9�@Źc�St&ĭ �V�k�3�y��L?�p@+��w�l��[z�3���8&�G��$��h�v���F	. 
���.f�&��4���9Oե%���$I�k/'��=��E)[*�yo�j��r��c��gogN��T�T�44�2j��j��i)}&:ee�)�� �e�w�|w�.Lv�I6�li
C�a���Lf%����J�mUhU#�*	��n���+ʘdu���z�f�U����!޹��&FY�#Ky/�L^�`<�I��!��T�<�现as$	��ɻ���P��JTX��8@wM�I
] ͹u$юl��*�C ,
#Z�m �5�|x;�L���@��$���I��$DCHlzarUE�����&���3�Ӥ����h1A��6|�� �^�	pȲ!
��;�>Y���p�ň�K^��a�N��̑�A�5��o7 7It�4�z�� [B`m'��[����8��-H�c���qp��@jM�v�0Oe~��U��&���N��ͲT��/�JgBЅͣ��BA�V9�Y�@�)+A ��⠌�^\� ���$~!#Z��� �)�]Y ���@,fs�!|�F��9JY��u��c���E;�
_�w$S�	���