BZh91AY&SYx.|� ߀Px����������`�a��  >�q�v� �T$Q4��&�bhiOPm i�@ �4�H�� �4    0`��`ѐ��&��4�jOE14��   �d1��44�h   h  "�@�S��OS'�3DbF@Ʀ�n�R^�
�@�*�
7�kV��6T�BȲH
֢F�=j�K�Z ��Sr"QJ�YO��ׇ���Q�G�~���������������������i
a�,$���K�=���ȗ�U��C@g4��Me�eZs��
�APK����W��4���/�ܒ�im��YAB��K��N��l��[*X���3,���IǓbe��P��ɬ�D]�%Ƹ0�*��46'��5��aI�h+�ՍSA�'(�UB4B���Ic=��ֻҠ�/��쮂�j�Q�U���J�i�D|0���澈y��Tr	���I����T�P�%���0e\�ܻ���J��w^/��R�SI@A:u�TZ�W�qr���r�%τ�"���}��x��T	�'|���@~��sZl_+�uA`�:�)�a3�Y��Ե�0�z�Xh)����]bVlkA��p+�h��P���q���GD�>�V_�5�8��O�e���k4���^�̭�^�S�^�\��cSS�s\�4���$��8�P<��a�4��u�Y*�i��.�*R�C�u�%fSX����0s��ۮ28y��3:�9�=���ҥ 1QcB�=�t���^�*B��8�K��p�pT�_6���iy|}u�8��H�P��Ǹ�uY������2��P��|i���^�(W��v��ѽ�v���M�$q�fFEVE����(ŪT�!�BE�DE�P�+�q8pb���Ȳ����Ij��kXՍO)u)��r�B��"I$�w�	���"�%/�Ե��c��Y�*�좈9�
$�@��Lm D	�	9�F,�bC�szו�'�HBBPiX��uRF����'�X�\�[Z��5��l���i m��d!{��=T��N�<XߵP|m���>���<�Тo:4'�ٗ�^6*�SdJh>��#P�p��.t��Gj��9Ce�.�<(�l��i�b	A���m��v1�%;O�:�pf]~e�9�u]��Bc���$+JX���M��G�6BP�=��/�>����fI����Mz4�v΃�VW�X}�i��)!, 0H#!� ��EK�l�TYCI
0�ۛ��
Vk�'�¹f���ETO��D"`!�B�Y�L�U�J��K|6�*�5B�M!����L�Qv	�!�@9�����-jܙ���(�\��d��5���3h$fQ5=U����t-Z�+3임�^ebHc������im����u��!�k�A�J����,&8r�7��m�s�r�%0,����� ��Θc�\dY��\f��� (�\k(�B�$]C
3� �{�!p�վ�9�f
�3�C�F�$V��ԍ��b��qߥ� ������L�p�k��c<��g�~`�
u�n!��:� �9+ł��:M�Ue�/��_ϛ#'p���)tA8p$,���if��g�r�qD�4JV�TbA�.|TK햦�ΗA/wDI�pP8i�=ua��Q���gD�]�����#�=�N@���֢~6-�ɼ�G�
cSw4�Z!=&�Sgek���l�q�[р����"�(H<>U�