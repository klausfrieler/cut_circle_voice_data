BZh91AY&SY��f �_�Px����������`�pvR�   �n���zz�Om6H���4��b���<�  h�@j)$�����  4 �S�M#&�# ���4A�e)� �h     ��z4#&��OQ�M  @4JAOD��S�4   Hz��fX�}
�����a@��_U����Y$A�+@�+?���UJq�GJ�g9N�v0�N�կ�:���1m��m��m���[m��m�-�ݖ�n[m�m�{��gw[n�nK��m����#<_�`|?�T��9������}���pm|��(�J�s�qp%*�tfDZ3[�#	�ʁ;�hX�.*�D����4x���.�p����ڮ@��/:�8l��M��"���Y<�JR�і�������ˆ��i3v�f�Vm،�u�W/�xN���:c��j弾		�rs0q�]�i\��r�j30�0i�f�*����\�D�Z�Ӆv�i�i�Z���g9����L
[���6<�ʨ�%��k����w3�h`�?o���EeR�g�&���D�֠��PAj$!����8��DUQ�E)1��-jI�Z�H�v � B|��v�cq��_�����=��A��rH��ޞ��
�!��<>#ODN���X���c�EM�l�j�';Z*WnL	+7x��x�M�lC���c��7
��Vf�蜘�]��T�J�y0�: ]�|���l멡Y�7�"��׾�����و��9��(2}ي<.�2�c��I�<�����+���y�Lc� Nvq	7|�?6�@yg�	0�����i���rt��\�[�9cˎ˼������������>�9���+k�{����+�ce��V]#��"��ԐdA����ϱ����	�" ��;�k���D�@�<�^��'�X8,���p��DeQ��r��b�������x,�Ȋ���K��(9O4�*�P���N��F=06�#7�$��Z7|ˑT�s�W����{�<cG�"]_j&hc�٧;���{��L�1j��d���QK`z5�|�T�*2<5k�mL/
Zj­@��û�y���E�#�Q3֩I ������VXwܪH��Ķ���3��t������d�FJ�E��B��9��
���-@�	\�m��3��nyR��\:�-��D��kPӝ�J�t����y\�\�2`=�|��Vp�NH��@S\$�*�	.��E�y�J��w�<�������n�H�����뒻+l�;�ZY����s�^᳾�e%r%IP�@�KH��˝<jwELT����j�`P�9������"� j�����n=��1���U�<+��R%`��f��}{�,xV���_���δ(f/S\މ)Q�H����ʅ|�����{|�����}����`,�G�[��}�Y��X.�C��
B��QA%5Bd
�H`���5<ۺ���{��9��Sp�B����܁9<�f�T�𡃯��BX�;"�<��2Mg�`Syn�p����~���rv_�3Նz�F�K�����`���x�<A��=��C>��w�9=��/ֶ��D�v��WC�^�Z$�6�-M�{P�ŷ��kîo�U��S]���a��P��<��y��N�GB�D�p��Sw}���l�=��Vz� V,�A��l�3S�^F�[���)��{��p{x
��C��{}༎��œ �9<�{�sҘ�]WV���>��BN0�@�+A��q��
��WC��d�������(cp��hX&���d�B���`��I.��^dBY���B� HX�Ɣ�YHR
��*Y#��P�M�%TD���vJ��EHe��aR#
FUX@ �Ў�L\$6�M
EBb¥Ūā!H� �����&���8�mt����"�#!�u�7�.n�n�xWG���)u2Wѡ����Z���M#g�D�X̟��B�	�y4�ۺ��1f8xT�S`T�%ܫ���j�����8PV�U�*X�@����/Z��7ظ�'��hPe�	)��TF*��\�'x��!d��}O<S������P�EB�"�x�=���"w�@ ��iwh���M]���v5���0HI H�@�(Ym II B$�d� �^��/C�
0��LC(VԷU(d�s��*jX|�AJ��30�I�ȴ�Vk��%�y�E9��@�ɳP�}Y��?kmńAZsh�W'R0�M���p�I޶�`J�sDE��5�d�P����6T�V�]n��$�22BI��ѿ�Sr�~����&)�z��I$���=k�&F��dr���u ��̺h��A[٧���v���@�݃�T,
3�JRH�?exC�g,�z�iY6Ȍ�a���e�����I����k��$lՉbBIT�y˲'B6pʵ���溳�'�22F��q�f�i��-�����/��Дn�rf�'ԳACH��M�	�	q�ga@�*�X��U�T:�Ś��*��B��e�L��ͦ4h�	(KF4�*4��=;�LC���[��pEw��T*}o)��H���;ʞ�T��������Y�V�gElJS�#�i���M<�() ّ��H��!O�rE8P���f