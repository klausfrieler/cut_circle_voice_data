BZh91AY&SY1��k S_�Py����������`�p��Y�j�5;j�� P �(�������@�M ��d�S�U?)��ꆞ��@4M�4U%0�I��Pi�@�6�0���IM �      $҈��S@C@ �   2�hz�d� �h ���  %S&�<M4�z��O�6�=OS�@4�m�Q�=����j� ^�U�D??+ W����1�BBD@nPR4"u���**`A��U2R�����?����>�����I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�$�$�J�)$��IL��������,8���w|��=��w��t����M�$k����E.�K���G(�̨I��d&��^5���ba�ݼ�$���0�t�&0 7��n��r	en�J[!	ۇ��0�`<=��
��O�Dkj�{���U�1E�Nsw*L�mAD0��rbi�� ���y�o��O2��!ɻ��Ҭ(�B��{���eCfm*��I�q�I�����a/c�b$C����2FCkg�]I��r�D�,m[L��ͫ���@�h^�N�8�r�d�+��6rqؼ���5UW�B�T��q�|.W#�rYZ�ʫ�T�HM�Ư21�	[Zt��	�1G@���� Z�����2�Zie'�CM�Z=3�jĬݫLx��v��j����P�[&"-f_���,1���ǸQ..�1��eF���E�ג�I\�XA|���������2Hd0�=��X�b���n�w����kZW ci���7����6�_�*�P��/���za�H$B	��o��P؂�����y��ʝ¥�59���*�b��^�i5P+r�̌*�)Q�7i���F|)ǥ-}^5�إi敋�5fy�d��ٷT���{^�������I|n��¶��LP�ljS�2kiҭ�jg������\́��,��ʙ��"طDyș�P��� #�}%H2�v�ָ@F�=� �� ;ѳ�AW��1��U����h����x�D���ٳ�S
�Rv@����T3�:�f�NY�r�uvf�c�8;0�'L��e7M�ښ�3.�[ ��5�6£���ߪ����]s����Gsѹ��h镁�r�y��,�U��I%���N�f4�HuD�!.�+��a#�s0�6%���a��lb2����>K{Sv+��;��J��C��WU}�W��m��7gS(n�c[��㛶�����a�E8~�i����yfs���/:���E���I��M�y55�^�z��lOH4�����WVۖD-P+&0CF�l�<�>9i��a�P/$]�>���}h���3�j�orI%�q��Q��?�Z��
FaS��m����o2$�-�&��P�}��o"�y���v�v�����j���(;�4^7��i�9�2#�9���9��K�+;���R�$�e���ci�]
s[k�:�v�
�-��Y��3D&V�����JkT���W/���$��چ��S�N�˚f���e����NZ�9f@�#����L�#��f}�qGQY�5^��Wl�a,݆���^v�f�<��|$d0��,�Lњ��;b�V�c�=���`�V�n)t�
�kzg2"�a�y�4H�%��-�L4�e�D.��]�$�[�a�æOb/����jŭ��vl�~�]Ζb̲-��Y��茪���U`<���>n�y��.�#��uv��q֑���B����kC���8�1l/)�>����7r�OYǗ�Kcaا ��E�D��b�mN-Z�I-ʆ�u��UMQ��lם���2�++x�$�l�[��:��Rۤ�s&o	ʥ��96�ɤ�e�|�����-�6|l�--��kڎ�ܰ"3a��9�7���m����#��~5Vo^����R�F+���1o�=a��=����]a���n���o6�y$�[3�q=n�����`v��-3���8bq��]`6ڣ�4&��-�W��!��;cDٙu�	�J߸�k�Sn��/�sm=&h��U]�,�k?ێ��Te��0}��"E˳]���dXT3!�� � �S���ո:�$!uC���D�MG�m��g,M�e�o$�Hc�E�)VK�&^�g|�y�Z��&��#ߋ�Bf���G�ŉ_/�
~1��(Y��NO��?�))F�dc��V��wg#^�@�y�y~m�S�JZ<�^j�q�9T�ܯ�Ƹ!�M1!���_����U�l���&+�'����x�������ԒIQ5���q�;F;��5V��6���|�/g)�"�!�����#c���Y)0���S}F0��'��V�n��H']�x�͌�����u�[����y��w��׃�O8�#�c��];�ǧwk��%�yY���C.w�����#����	$H�
�C���N���YAJ��t)!�<=C@�.(D:�(�Ι
S	�D��h�RڅaUm�ZX*�(�R���ȱ*QKh(�KKJ��A�w1B�$pڒ�(�m���d��l���J�Jؒ�
։R�wb�K]�
b�ڥjV��R�(4����l-�iQ��h���j[J6����УPӄ0֥JV���(,�PFV�T�k[�	!��/IAKl&l��$���Pq�L��-ra�<K��|A$̐�1f�6~0��?9Ze6�t�������O��P���m���7�����-�ըN�N'����3��ƸR� �D ,�ŢU�G���K E1S�w�!@�	؞&�?�`�	�(���Ψ���M��g^��/ԚaϤ���ia�SlGa�E��͊�+���y���z� BR�E9�	-�5\�ٞY�9�o��v��"�U`��V,P"�[aTdTb��#A�"�V#	4!e��@0mOF�v���n{�<�x\c�;�%L[��EYj2HAIS��d�t�a�ð���PMٶ���x\�/PS���n�����XJt4O*p�܎d�a��Ho��Gڻ�BH�vH���#�9�s�a�؎�Cr�߳�M���$$0�<[��M�p�V-Uэ��� ��FI	"��=~��&\9^;�(
�C�fPR����/-S%�5��/T�Y��dF0� [��þf���H 4�*�!��죳 � ���;�4��.{��T��%���8�:t��'���w,�`$�<�t�X<U��2�<������i�݁>p���H�p8���"�q ��p�O:����5��|Ne��b��T�4M�i	�\���-�l�6�A�u��xX����Rܦ�r���d�"��,h#3e�����0L9il�Z����K�T,8��L�S6��O��S�
�C�>;���)��t)��uv���66�?�6��J#�N�2����"�(H�{5�