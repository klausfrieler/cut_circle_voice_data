BZh91AY&SY�R�� ߀Px����������`�_uD 
L�Ƣ6�0$�2��&ɤ�S��� h��S�	���h�@dh   s F	�0M`�Ls F	�0M`�L6�O���4�3Q�   ��DAh���ɓʞ��C@hh�mCjSI<6$�]BEB��!n)@�Ԙ6�I eƗ��}D@�	���M��9ʖ]\�]��k�gGL��<�B��(�1���l��=�L3�n��밦����	ri�]�іO�w�S� g3e)�B�!��dSS����:|���[u�= �4+�ٮ�������x"����Q�}�c�
|#Pnfr %r�H$r#���c�Y�]����6Z/��<V��$���Æ�K+�50�lܢ����J�vJ$��6�fY��q��fgl̉�]��7���`D$��!×͉m9�br�G�+�hp�V�I(G�s&R(C(�dpCOB�v�uvx�aEV���#Rzv��vK�6�J��1�(�<pa�L�=<�^܇��An�C[�v�E�.䓘��y�Mo.j[k,2a���W���kF��6uA���wx`�ڷ~���lޚ5
�۹L�Fj7[m����Ƃ�b�p$��A���:9*{��̩��f�~�*C��r��5f؄Ǐp�+�k��Fš&w,盘�!�w�M:�s3#���Fp�y�ӂ��a	,	���lq���T����z9z�e���<O�J����e��r��i������m�`{�+�9��s:{ֵ����N�=�`�%�dtN�w!2�!; Ő+AR($��1$H"a]F1#m��2�p8P����-A�e ���?���eqg�h��Ѣ�X�g�b0 �E���'yi��,��l�;j��CQ���|h��I�F��Bd�zw7�6�F�y	���3��-U|�4 =�fx0_`T`����I�pm��w���N�Z�#�vցL�v�'�����Ey�p6ڈ�HYpU�W�C	^��FL.[���q��Q��"��լ�^��9���5�*P,�[.�<���BEƐS�$�H!1�8�.ɤS��.�5��$ȢIrHL�����C�Lf)�Ob�%h7=ZrȀ����Ixܯv�3���S��=st#�Uf�L6��ܗLV$�����+��'�=1�!��T�5�OU�JÙ�AŻ��P���'*ǭg������f��&Di�@t���Ie�vi%8F � Z0�Q�O��Ȫer�39HF��W�A@�@�&DCBm���d
����5��4�(5C�LŪz���@͕6a�d�����Ġ�g�X�Ѱ��m6t����Ga����� 1�%֘���E�%
��1ڧ��J��	lt���Ӓ׬pH�i��{�{'��Mժ�z(��y�POx�2�IQ<��yYz�r��q" �ג5͔��6��!Qe�Q|{��OHI�`�nI/��yJ��[�hss��[G���=��ٜ�8��HϷh���ܑN$2T�q�