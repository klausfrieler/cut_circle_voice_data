BZh91AY&SY@&9- C߀Px����������`�Q��      
 � .������MP&��   i��
h�m��!�4�	��� �`�2��I��I� �H�   !��`�1 �&	�!��L��R&�4	��L�5M<ML�SCF�M6$�K�E=���X*��)��Ԭ���7�
B�D�R���8�/�H����d)\���4a��ݿ����[��      ��
�DB���1P1�     � �H���(�`` """ 1��U�)��>F��sۨ���7��&��}^��5��T�!n�rrK�21T��Ŏ'-����R�De�S������"�z2p�3)�����y'b�2u�`H;���B7*�䋁�oP�!c���W�r2wT�×#]@�FFM�T��D�[�[Ծ�XʵN�VFE�����m��cj�_T��b�o��-��9'�|�������zMW9Uܙ�y�m���ԝow�vW�b�DN���ASPE���i�t	5;FƋǀ��9�Bʪdf%D�A��шS�8rJ������.S��F#yU/]�A)Ž�C4LA�+p�Ο���c�F���5�ђA�7�b�U��2�w0Q�� �bۥ��ma�vi�c�CmӬ��n\V1F�I�y��pۏ4�-��.����̉D�q��H  ���k!1b�L�ƻ�p�Ĕ6-�IU����-Iޖ�g���'�~��u��ӹO�e\-�������%��V[��4b�_f� _�.]���h�R��I����V���6�2�B�	�p$;�.��#9T	$Iَ*h��Kl	5\�
�f�����܈��y\�6��&��Xk�tA�^P���u[p�q�1��!��ǈ�vu��3���ö����cl���	 e�	�/�2 �z2Xq�����m\����j����ܑ����
`h�A8$!,��ؐ#]���gT7�&�QT�e����e�,��3��/OШ��)�x>�&/��Ou�" �_U���������2�sB���͒!nX��@}�������YU��zd{<M1aN�?���e�9x��N�6�-�&^��bq$�@˟@^�kN�t�#��I}��TP�i,�S99�dX�zo }-�hI�)�@��XI�<�!���&���ǝQo���-�}Tp�<���&��n�Cifi \�{�}���}5Q���t2+������bm�KNd�Cc��T$��f�vz������L�A-a���=m���m����Or��� E;��3A`j�a�L�' �]ş`t|��@ ��1���#�0��`��>*���5;�$\��?yt
�S���iQ�4��5�*�1#i���"x;�8[���!G�����}���2'ޢpE��TMK�D��|'r#���v0X��)��E�)g����7����\��̻�#(�w>�@zE0������Df><����,ٔ�����y,,���U�́XT�6�#�R8޸�ͳ[���=�f�Q�f��ZP򱆈�A2��%�膩`�(Tל$-�����wwt��u��Ve�ר�겧׺g�[6����Ǭ9)B%�/�-��3�y�3G��u�:��������B��	�Fq,�vf�Gaށ u+��s�������q�s���|z���\;뜨�x�q�`��]�x�r�=���ݬ��]xE^F[�YEec�C����ƣ:oj�$�Gb���jdl�m�M��Ҭ@D�n�;�~�c̹��#����#����XLk([��4Q��3<\�Nk�;V0;#�^��n+=9*#8Uazl2@��+$@��Z�*��=����F�+T��"��M'őR.���B1(bt�D�t	kq+u	��`S��D����Q_'�A���s�wѽ�2�z_�{d��_]a
0��}d�����v������rf�1�#�z�~�u�վ��wuS×땑�er�O!�D�C-����N@��YVm;�VL����Һ�ft�����h�W,��GE�t����5ן�gαF*@�I�
VT������<la;��H+�OD�G �[zȾ3�No������UG>��34�Qi�؎�t�sH�;)���8C�������m�{o�����G����s��۽�:"6�Є���$IW9&ӈӘ�S�Qw��Iw���bbv�cp(Uփ݁�w̞Z�{3�{_�\�ⴹ�;��}A�O�DD@@��$yt=f�olx�AvN�Ғ���t3�.��.XdCf����Km�0f�2b�(�VVTX6�TP�Eb�XR���1�R�[RQ��#����
��%b([AaRH�eI+ ]��E���
¢2�*IR,����L2a(�QZX�kX���.nb�"6е+mJZ�,X�,X)R�ڛc�k+�W�,RѰT�n�ޛp'��a����+!�}��@!��o���O	{-����w��<ru����5�?_%�ѕ��γɼW^�_!�$][+���3���l�iō�"|v��Z���>�DK�D�V �qf���CF����$�?��%�k�7���� �nt�������$�p���o��2p����~�wr���i��]`B��&ql�\i�3��q뿥��0&��H��F��X
Ab���
@X
�FE ���EH���VUXl0��h�`ҝH#��l���F��l��?�3�0!��"�T�A�"2�q��n���z�c}��#����H,jf ��aN��Ƭ2�@���dD�N��M�,�Z���U�znwL��&��Ӱ�����5��%��s߯��D�r@(�E��zhc�>�]i��@H6� R|�"w�	u�l�)����Ă$�(����"R�Y!�<"������buu?s2pn�m`E� z,����36ڜ�ʙ�9t�nw@��i�u�F���H��T�����a9����x�"n�5o3NQ��_-�w$)�����y�s��D��w�B��M�"g
�D�C���Yˊ��P�=�r%qP`��$�ڢ�/9�.h6��N�88Y4��e)����G5��܂%��)8��9�d�8�E�a0��ve-�D�RvH�Po렘}c$$��c�3�&em�3 ��L��"c��"%����"�4�+ߌ�R�=
a٘o��ܑN$	�K@