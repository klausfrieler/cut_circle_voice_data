BZh91AY&SY�J�] �߀Px����������`�Xp��s	u��T ^�"AT=� ���j�l$�
d�`��z�T=5  � ��ER��10 �������	��S�M��h �L  	4�'�      @��T���ȁ���b0`&�F��@��x�)��1���Ѡ���Y4U#�(�5*(�Pp��5j��J�H)"�T�PG��f���#��Q� ����q�����.<����Z�n����ԒI$�I$�I-J���s7u$�I$�I$�I$�I$�3373Vff�fjI$�I$�I �I$�E$�KK330fbQ�� �!�y��q�~y�������g���9��m�o�FŬ˥A�neaɩ����,��M���L3'��n��uP���0�Ҋ(N1".�ȓ�n&kQJ�-@�w<G�1��ک��Up���x+T1"�f�:�Qcy2��(��#732��g��b�n��N��1e⫻�ڸݙJuN�\�2X�W�d\��ۗ���~��?�(Q[=F: ��r'9̦fᨦSg}mxॸ��L͌#�U���Z����W�(L�V���ŹGilırF�bT�g&���w���B�Bj���N��33A4��3�`L�V4��1��� s���0�4����<���k�<�B#��&�Nk=	�MoX�7�p�9"��HÌ�y+j�[�/jd�S���-�Nރ;U�v���,Sn#vjA����6Pd)�츬NC���םy,h�Ȯ���ڴ�3�m���oA���+�̡�C����<T�<�E=�K�[�А����V��9�|:g����}T�玬�*�0�ØAx��i=��pE�֡NpnJgg�DS������漩�!ò0���h���wDؗ�A>�}�	K�����n��73u$�7wc�բ�����&����������_a���BD��%E��{|DP�A#� �ު������x�L*��M�%/��vR�H���ّ0_. �e+��]���F4�<B��z6'����\4��@%�T���10^5�#\�l��sm�88I��b+�ݍ��8B�m�<�G��v�W1�Cp68��C;�aino�7�L��Jn!��=|6���>���Y`�{%t��3R[��`�]]�Ӑ�`�|������mL��)�)R�� mDP���%k�������\#�BDa�LNZ�,����A/`Q�'�qg��=x��8:�X�������'��M�xDz����P|fC��6����q�:l��Ҥ�滴]]V�id�m��85i�PnƂ�� �OOcg����K�a1��{)%ڷ�I$��v�ʊ��f&ȗ6�q:�J�Fa@�R�F�p�)P����{vi�������s��k[�)c��> b<����EZw"{��P�Ǳ���W7T� �GDf��oY�_n�z8�P����0�E�G�F� �i��R���YVJ�yB��#4���]�A���/lo���	$�K��,�d�"�eC��OW-s����KB���(�AY*Wvh9�e�/	�ݢ�>Pt
U��/�@�;3pK;�lǷPW������H����o���8	��{:r;��L]WcY�Cn�����D��<����3�<������b�٦�M�c7C�iDÊN�f��Y�qX���vub������޵�x�w�J��q�K�.F����B�x�����T��e>=�8X�vt�u�
j0��c�J�3�û��}73Tr�W3a�iO}<_�Z�jg�?s�n�w]��5eE?����'5��:�`��x�1p�"ī�g'�H(��C�н�覡��)nfb��*�a�t�n_P&���6�*e��ӽE4�4��4a;A��-�2z�f� �n��4������k֋l:n�v�dk�{ih�ح�}�v�W�;E&����$�P��"�I�Jt��m���YM�/���@�5�o5[K�p��NL�<��˒I,��;5�B��@׃f�DC���7��M�-r�E�1HD!�H��Mt�T5AT��#B�":���	~{0g=P�Q*����2����ȸf�������R�+�`�{��vZ��������I�|��v����2�YbM<���g��i�!�3�`^��f�3330$0�njf��8�<���0��[Uf#�.r@D�����^�7�ť��a�5UC䟀��0�
��O:UXq܍c�:�N����A�N�(d?��~1+5��_���Y��f]WB# ���2�Ub>2����Ӣ���R�~�R���>�1��Ӹ�W�11�ܳ39%Vf)�y����LL������Wj���I�kZܢU���P��XZ�&�7+I\Pe��j ��0.�B���<�
�t�ֻ����y�0�;��P���4wl�:��Vȶ>7�'rX�]�\A���>���3u����1L��6��*��hMl���}��I	?,��!$AW
��+���2�D�6��(Q���'8��5��LJ�ڦx�cS'qj�Z�kرJ���E�(��eh�,V�Z��D"*�=���ɵ��c+,`�	[�-�P�2ҫ+
�eb�+$�Q�F����+%F�E��i(#Z�FJ����ۈ,SZж��J�[b�
�*-HԶ��L\e��,YZ�(�ʅh�PZ2�ZҢ�b�e�]�D�T�j�͔�ɦ���(lf��ڎ���$&d�ř]�&���z��V�_��������j{O(Z�_r��E�N)�h}��h��	��~ߎ�Tb���i�Ǹ�EN���n��ôv�T�UOљb	�b3���j[�@�b�����Ne����F�exPT���X��iF�5����ҕ��K]��'}�}��т�R��$xߦ��F�Д]F!5�w�� `KAk%F
��EFAb��Q�b��H��X�,b(d�*DPPX��eDBI�NJ@�Ν#�
蚦2�w �˂�b�<D�@�6���m�I�N��i'�^�ƒނY/�- ��l
�ڂ�4VS~��;n`�%��m�9=��.K:�F�j#��v\�#�v��:�5�U��hw��.���	##��$�����u���U�S�r�@��� (o@�=�W�&E�ҁ���T	��@�H�I"��X���Z(�����*�\,�P�ZA��+�A@�@�%�DC�b =зl�ª��ڙ;�1�ɥ*�(�$4X���jF�ɍH˶ML���1U-�A�p�a>�c8�%�F��D��vm��0v�G�������{BB*a�\���*
��h*c����.�c���-���ҋ6:����*������
��׊ƐE.n��SP�����I_��;�oY���\�@8�lc�V���2%7A!Qa⨌��wZ���Oa'I����O�
clkSNA0��ד���O��J�?����n���F^�"��rE8P��J�]