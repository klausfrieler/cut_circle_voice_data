BZh91AY&SY��%� �_�Px����������`�,E�     � �1����S�4�Ѥ 4����)�`�!�L2hр�&@� �`�2��I�J���`b  	�C�0L@0	�h�h`ba���A2i��ɩ�Si�����أ�0�	���
8������k��j�p�Y$B�P#H����\� ��#���	'*���gk���r�'+�s�Nf[���ff>fffffa���̼������Y���Y�����333330ffffff�������̬ŘNfc�NB5��	?D��_	����/-#�$"���f
]�R`M?�دKDS��uj�:iv����t����4L���/�V��$�D(2��lC�=� )���{��3)˙"�Y1p�Usq��S]�����4�.q���SI��	3+2�Z�e����#0J�;(�zٛY�bD�6�cJ���7Ō3�8�����1�QxW�beV;]�����kf�>2���S'"�`���t�%�21���fY[K�� �a�Ř+���p��S3�|D�J�HЏ/^l��c�P��u:xhs����9g���2��o�X�L�3@�D� �(T\p�L�+/��
����r��3P�y��|���  ~�,���r��7߃����cd\���I��zU�Y����H�ئ�3[g���(�8>�珉�~)�epw(�L}{������4��F�	z�|�WV�'q�3QP��9��M�f�?�q9��/wݽ���ilR�Cׅ�(���Vǯ>�<!�ƞ�7uu mc��+�D� qD~�2�"8� ]����Q�N�C�V]������
d�k'ni����`���DKu4��HD;venhe!F�	ǎ��K%��Fl����ɔ�MI��i�٘��lQ��gz�7�����S��4��婆^0Mv���M�x�ҁa�����όy/�	����3����@k��wW'd�6a�	�Vc^3���焊���!G�������X��.��� �d�9��cM�0����F\(��|�����f����l7J9ɉ�}�Ov�g�O�L�0}�}mX�]���Z*H��ʘ7�c�2����ʄ́lz��y}�Ӊ�C'�M]$���b���m �U���ܟc����
Ǡ�T�l�c `3NAIT����v��7ѻl֩�c�I���YtzĚ�s8S����Q�_k;�{u*Ŭ��jӳ��plhul�� �;`J������jN�SI�	㏶@�yOt���l���>��`�±z�D���G>ך]�	�uk�A<· �WKvm`
<����{�Y$Xs!)i������[��:���9�cr���3wW�^��˪n��QX+��cUJ�����	�=z�Z��iJ��<i�}���$���[4Vdr^I�Q�@�]�_Î��cUY�l������mBZ��|tBB5�\�
uT�g�Q0񗻝��i͉Q�n͸���ށ@�����h�(�ă�m>��W)�b9�W�H�Ws �&�E%��e��h���#�n�l��]@dE7���b�ES�*`6���Ģ�s䙂��@Am0�m�v�0ݛn�&�z��wa2�r�)M	�S�w1� ��
�H�O���֍�M���;�j�KOe�벩�\�n�=}ۖ�T-�BmxU��m�o�ozu��ɹʐ&g{:r�3�ud�MD��n�սc�#m�S+٤18���F��[��`"H"M�Q�u8'���&L��)�P��M�ǝ��
�O1�'�˦ݩ�B�]sXǫ-�ļ�iع~�M���l���|��F3�gff�2;�c0қ,j�g�w�l�x�NH�>1�q/<����w�@<1QD��Tw5��W�ja�����0�e�C�{�B��)��T��Ⱥ���d�u����K�a2y��# �q����G�$~hI AP(P��>�g+���@���[Z�2�:���AMs�V�e0ª����ҵ%Y"�[BV�n �6�F+++�A���R�kAP���R�XE�Qa[���*صR�km����F�AJ؊��V�)�1eA-��(�J�-�KlV�F*�82��0�i��-�-1bɌ�T��5(�*[B�����rm�>�f3W��Q��&� �&a�Z���C������Ƥ|3K;S����D5�����rM�Cݽ�|�OBv�9}Z#Q��S���&�^$��XW-��}W��P���` ��mY
 �o�o��7}���R��?l�tQ�ͯ���pگj(�N(x�I!rRɞ�Ȧ���W���+G���蔧}��`P���愀�wBޣlh�()H&�N�\1��dQB#"�1"�(��+*Ȁ"�PQ�X�,b�Yl C���&)����|+u.����v_��Ƞz*$�Ց�B"����M,5��g{�HOV]����^��/E��ݚF�ٸ�AP)��;�V�*6ݵfѥHo�.Ź���e7����.4�6�>	��7�Wi�^���@�q�!/>�筝�J�kɓ���N��s`�}h�}��ŉ��l�]LN�2��\e� :
h*�i�3�L��a�!��(h1;�����7�mI���f�5&�3m�Ќ��Ñ��L&��А0�l�I��5"�9���߷C�Aՠz?�r���2�m��g�VZ�j7@o2G1���y�n

��w���ޜȠj�@�c��Ŀ՗`����	�BXa�q@�*�����cJ,���z��E,k���j1 ��.�����Fy�`Ai��X�D8�{�Z�I��o�P���&^8�T��%O`T�q�4���mN�g��*K���|�i�5����tR��^�����"�(Ho�� 