BZh91AY&SYk��� l_�Px����������`�{�v��r�B[Gy}�;���!$����0�=)�zM��'��h�����$�1�� 4�M  �F�)�      ����A@F��  4� m*S�d�D6���h�!��H�FQ�4M)�oQ��4� 1-$�>��$@�P@�K��I(�:gԘdU � �C�g�'�!4!�u� j���^�h{]�������I$�I$��RI$�ffW��$1Zo�����L���ݮ3�(����M/�^�d�c-J��(S�f e^�
c��������墦�'��V_�m�g��$�M&`SF�6<^%�����z��q(&�P����e���v��R�yb���,�@
_J�7����Z�aPvV����A�d�(*^YQ2�3��\[�$1�r�w*�`T3R|���AE���V�[9��R`��u��̲�M�xDlƢ� ���j:��s��o!��<�VFSk��6�u;R��4�9�/}�G6��dF��wc��r"�Q,+MoBa���ӈ�m��gvi�&La$��Y��gܶ�0��Ϳ{@1Z�m�/N�D��4�dD�7R8�C���2d�Ls��f�Y�͌7+��J���+
N�����3���P�n��Xк8v����!�Q<�'&�m٘V�d�9�6��ص�\��0gqǑ��5|�I��n7"�Wd�Q��D^�qa�9ȝ6ٛ�Ɍ�5/�*"�tHZ�	�|�aCPSi�r��	�J�7.��KX��	&�^M�	P�Ȗ �ju���eh��;z�c7\�%���q-!�N��״��6�p9����^,m��;�.7�#p��7!�*:�@�
�G:�>�BJ��h�N-�ڱVLaFЅ�lFLkD��P]�hi=��R�i+3�,�¸����s�m���C۶���60��<C�H �^Z*�(��~p��W�^If��œ?�⑧x��k;3I��T��,V�a1���ٺ"��5AMSbЖK^剢��5�(�!�҉�3����Q�h��Y�F�$�l�V�0x��羞2����ʺ����G���>i#��S̭�0M��o�k'SD�;̐;���Q�+�'ؔ�.�T���ʹ��|E��!}͉6@9s�?�aʞ��u��6$��1����
}1p��V�C�EO0d��L��މ�<{+�����0(@��K�(�G5�7�����
R
)�;l��!PX*��"�VD���B�(ށQl��R׫����B��ON�b	��&l�L&�[�ԋvii�H�[S�δ��Fb�pEA<"�G�$�[��´��N�վ$c&+5��p����*đrL#;t_���=kr���e.�k9��tt$�Qk���&�@���4�(�z�K�$��ڹRh��e��������H���PX�v �%Z|�;L�����\T4�A �@t�|HBM�G<� ���������6�c�&��d�n���5գ2I�y��򬠅K����'c8eR�F��Q^}���F��.��Ә	���7�� �J0$�ݯJ��F
d�z�E�ͻH�*NC��0�͊-_��U1z#9�I(Y�9�M>��H�����MJ���!�疂��`N7@�LV�LF~��SC ]��D�M
�#JI	��VW ,"� *��p�t�m���'s=�_6p���"���7�]��BA��