BZh91AY&SYH��W �_�Px����������`����E��ACM E	RB�� ��B25�HI"a�	i=4j2�  ��i���4��#F��4�Ѡ���J� &L   �� �I	2�h 44`#@ �0L@0	�h�h`ba��4#�&�4I��� �MC�=f� )=��j��` p=�+��������d�UK�D� |k?��.A�EN�AE/��ߑ��OGOW^����Ͷ�m��m���M�-��6�m����I"�H��I-ѻ�����I$���ۦ�v�m�m��-��6���I$�q�� C"�?������_'������q\��&��"��9�6��RTtex��M��YWQQ��qd��؍L��rn�%)�Q�cdM�EA�
���17�Dd�s��mla�E�8���«�۞!���ڴ-Z!T,oe���uo\�VDZ�������9��W16uyDʺUn6��B-m6(�
�^�P���E�������00R�Q[������hCQ���U$x����{��5��㗕
Jy�qG%��n�{.��ӕR���YC-sV]Z��RF��B��ʘ�A-{ih�VO��T۩w�V}�>��8.�D���'���H�/��)�g	�Dj��0�ZG幷�W��5-�"Cځ+%��#n��E+J�m8�6h^��f��J:�B兂(1��ʡ[.kA�p�
�֯��pqa���r�rʐE��Y�W�s����v�*���<����M�l�#�ذD�gX��	��蚩����w�C�_/�B�&��0K˩t'<.��)��YT� )$uN�[�\o�wL�ٹ�6jg,�okh�XL6��CI���ڎD�,,2�5K"���������T��{��z��͠H�읣+�E�00T��"݇0�/�ev";���� �bz��@%(��u3����\��f���ra˕���b�� FF��&!���M��@���:z��A����3����h�}ڏ5���l�pA���<���g�q�z�<����O�\@W-O:L@�u�&�o�|+�F��́xc0Ʌ[��ġ�������kZ�;�rqX��*��d[�t�j�!ށ0�Mb-��x�d�[+ 
md� y@��~`p��Y��D�0�A�À�ƀ�O��������h��˕5��!�{��F�+���ű7�� �W=��#�Q��@��"8H��"g��B�]:�� _#�3sk��	�a�r8)�6������Vmv�wz�D�͞6{��T��lT�^@���ٞ�{5FƐe7bMbh.W�|Jiې�x/�,G�M�'��r���Q�tB��s���`�ǀ2 ^�V��*x�����V�QC1Za�W��09
�x�#'�^�k@fw�=�ع5��T�<�Q"�*�����2hA���΋�ΡRGoZUv@!������"����w���Е�����kb5Q�w[u���*��p�<�E�W|fo�J���?HL�	�.�A'9p��/��@ڌ"�_*�@�GO �7i�y |x�������<�����#�����@������#7k�������@LH�أ���rO{�#��{G�
�ʛz�w��{�ߢ	y�4��Y�W���=%�[3�q��`v3[Q�5&�e����S�U�-QZ�,磠���kf�����BB&>nY �t߅�����{;�5�du���7q��!�w�&JS�bZm�7U�`�� Bޜ�r�M����/�R�w�ԒJ��6�3N�c����&]%��Fc�Zo*�(�ݼ��t��dY1{��'{��2&[���vEG�;�82{�b\C`͑��w���yD�0,D�ב�QELQצ��o����t��E�]��t��&2��:(�گ9�2Aѳg�ވ��:��>��D� 3����~�{�v�����9���,w�$%�)���"[2�lR|�x;W)�(�1x#��na4ҽK�iB��岪���R�P����Jg���.���n�R�
u�dǡ	���a���b ���6���ˈ�b�Kwz��M�٪�#qܓ�-̀h��^d��ݔy�u�pr9����H���>FEE�Z�k��(1�z̶Mc�ɫr�5����Ժ�ظ2؛�5��U��U}L�āW]�x2�{WӭM- �*y�C��=� �mDV�I���Vu�wͶ���0��}V�̫r���$����SY���%�[�%�\3��c�Q#����	��[x����v��p�q���,%&��]��?dE�1u�n��W/w������&��ﰃ�D�n^G�*9�"܅J��s��[�8�S�L�5�G�w�~S�QW�EP��P����y�n�,�%p����qt��vv�3L+YSM�Z,X)P�U�T)YX�(���Z�o�I�:rҨ*�+UmcdPU�TX�T�XVVBV��6��FH�q�9E�
@�6�,��B�Z����#��9j��E[K(�DA��k+2�]Ra��5
ږ�ֵe�((���Z����ˋ��Z��[[ye�m��[�1�mSV��Z�y�8����ɚ7�1/#���:"��$�;+B6}0��}��ݭY�,}�����}:b�ކ�6����:����z�I�}��Ѩƭ)�R�.�7�D�<����?p;��=��b ���Y
�5S��8��l��(���Ҡ��F�y�)ǌ��W�L2Nx��!rRɪ����>�L��Js!�u��W���q�����M����Ƿ[�	�+k��p^�ߎ�Z�A����1X�QE�,��1T�P�b�)X��B*,�DX,�Ȁ"*0�I!�I� �j{p,G].��f����S��>���L1.E䈲 �da$"�5���Ɇ�?����\�r��8����y`[א���O*%64®Τ�C�_q=\FK�됒4���n~��i��c����ӎ�<�؄�do�CC��޲n����;��b��ˈ(�()^dQ=��bg�ۀn��qT��;CB(��Y3��Pt�Q-sN����-��AS� U�Ȫ���X[RIk=��nNSS�)ٌ���Ne��1�(��f6�`���Mh�6�c��sY�1�����P�4Y.A�V��Q��˘��)����I�s�Dϊ�,"����Mar(��}~~&�11v�p����K�%����t���է475�'��"�X�)]MF$���t$"����bq,�.���C�7�
ՒHFD�H	
���TѲ$���N����d�'�b��\D�W`���6�Q�O��-�(|3��99a [�/Ϡ��rE8P�H��W