BZh91AY&SY�\�{ _�Px����������`�0��  T3�-#f$T�Й�����F�P�4�����5<�D�� i��    s F	�0M`�L$(L��FF�@�  0`��`ѐ��&��)S��MOSi�b ���[H�Ҩ+r#��b�����)��"C(������9��hJZ��W�;ǯ������7���fffffffffffff`��p��/ܰ��/��{u���ݑ}<�fal(Wb���F0Z:���77%�1����Sp��F��Ӭ��s_Ϥ[Ӵ��$VP���y+��[	��B�WH��)ME]�R�lr�騫v����ǐjGx��$ 'l+�$b�n�����T#ng\IBP͞z-/2y����uo��Z�c?���j�ƹTY��X�`و��VZ�Z��ǐu�g\L�V�4��u����i1�����L{d?g��L��
��
m�~������N� bd��� ,N�Am9 ����Qּ��?Mf�:���-��G�#�����h�H��̀0]�dΐ�!�N�	���la����GHYc����p��0�)���q�o1B�!�l�a�&QJ��"���<�d۩t�t���+V���,����lICk�ü2A�T��X��KX���<�DF���#2�>sN9cF�K��G,��[�v���w��4�l�kV�|i=ty�8�:p
��m7�$c�D���㍶Z���-�w����(��f�Α���~(C!Sj ����9hCU�[�ߖ��/��<Y�8�8ߒ���X��Ǥx�v�1����6c�T�6���`..+vp��m����ˉ�"ؒ�+�E�jҠ�L�ڡO��{��c{,m�i�:8�t��]�pr44�Z!8s�w݃��g.阇fe�BZ��H(�o[AFrI#lr*ҍ����A��j1Ѹ(�F��i���q*Ғ) ����_6tڨ�Wz�.5�5�,HCfmh�[���W�,�r�
'�4p�s����l�j����)��{��6��l��\N��a`�h��Kzy�#�af�@�_b��`|Gj�US�q�A �͑�{�4u�#�t�$��U�r�z�|��\"tF�~�6�TK#]֑�<�*/ƙ���s��r}��!-k�^�ͣ�im��Z�V�u�}jWc0m�
4���[�,�(Z�1�L�0�VW~�`+�J��(h*!�@�4��įv�&bY���*�f�jH-lf��v���0}�ŕ�Igd�uK%�J#ߤ�b�dI+�F��մ��@�@�Z;��f[���;��!M	s9��J|0���}�80��] �f���ѭ�XK��hqĤ&`j��;�%��$8�D���C��J0R�3r�LbhX;�ʄ��6�^�����Uc�MFF(�cNPe��b��yM!�ЌD!��H�ݝgI"�T�%�93���d#_HT�q�xx�#��M����!�$�_Uv0B��M"&�X"oP�vu�a�W�o��9A5�$	�E�T�9j���;�;��V�-�����g2Q���^"[J�bf#S����$T�y/�fR��RvȘPk�A1v��w1���	�[�L�'��7������Q/���R딛G��Jl�|��g%U�"���g�]��BBr1�