BZh91AY&SY�I�� �_�Py����������`
.�}*@  ��#T҅!�LMLh�#�&��4�����F�F��jy I*5=CA��     �&M4�dd�т0�F� I���� �  hd   8ɓM0�14`� Ѧ $���OQ�e?Q�=5���Ld�!�`iAJ�����R�����ˠ|�T@���!P���pT+!�p��)�&�p�.#W����������L����������l������wwv�w���������!\_��'s��{��O���ѷ��}��<�1��P2V�A��R��Q��V�qu�ь�� �KN�+��[S�&��(2m\[ٚ��vhu�Z�0��m��|9trU*�����2��)`miٞ�\p}��lڦ�X���"�oK<�\�vj�����Sp�!���=�[p B�5$!-�(>���͟	hD1�xJv���SB�~"���4�A�UYj"�C���z��;�֯�#q���c�*�2��Sh@V���w��/"QZF�)��Ti�/�}��.���eJ>�T����T犔@�w��&Z����Lݾ�������٦�� �Ktq�VG���#_�ܓ����p�����C�G&w'�i A1�b:�߂�qk����)K�C�m۽f#�q8�8sӦ����������C3k��4O�}8O��0j`-C�'���n^�5Q�d��d�T3f�%��8)幱�M�(rχ����b��%3���c*Z�$�'�	nw��ڌ�0�w;)u�WO�����B^>�c�����2�4�T�m�5������A�S�#dwĵ�����Lu� �#��{�<���|��L DH1/)3��Psh4� �q�RLz�R��� k���F㺮�V�U�����U"�̧�U��l���*�Ha�$B�|L���{J&�>�Dv"�1�g�*�s�:K�g��n��cY��*]B�r�aC����nf�,롡D ��Y�h:�f�g\*�U��H�z��T�j�N�u�{,��1ֶ��5��:������x{.�!�>a�Iu��c�]�Zq���QtPd(�>׫D����+�����eTuƪ�p"H�k�v ���[�-`"�Ӌ޸p6���������$�D���A�n�G*{=T��q�h��a��?ºՕ/)�󡱱���,m�4  ���>sq�tj�g���s���*�&��8ND�%Y�bLI�c ��ń�eB��+R�o�.�\�TXɴ���&&�-�[Dմ�V�2��-Kh����ʃJ�)X���EUDTTJ�m4W�V�-e6">%�,�Z��%�K��<�.MQ�?��І�e�Dhz>�ﺽ��o>��pM{0��rz�Wӳl�g���R	��L�N'٣����M����?WMō�����[����" uZ��O�;U�N�T��!�s�H0�9�����$���h<#���7�����cH�0�u6�h���F�4 u{Ji���
d�m�zy��m�M�DJV˺�~�.����ʎcD�]�Ï��MU�6&��F1a��H�$6���Vk#��1��E�Y��8A�2��CW߬a�4�!�b* ��*HW9ʜM��5��
d��j���|�!\���qO�Ԑ��疔ƄlP�d�gb5Q�;��ih ��'��`rjZ�፜�K9ę����ގ��#���W�y͌w�׵3�]�/����^0����$�.�'b�Ն%�%$�0R�0@���^w� 4H���Z|�^!D�cT�Ȓ@� �A�P�I#u���H�J"i	z�mT��𒵈7�����eø� ���B{��X �� A�#h�ZM �tolό�5����6Ɛ���R���]��p��iᮜ��ph�g�rbMb9tF�@P&t>��{�x��s�7 �����U��k��IM�	A��I�n���m![1�
�R!�6��v�ڴg�u���B�C��!yjܓ\UT*R��H�(['��fhH�i�:� �0 ��Ц��Y���|�3w���m��������<�\���*��ܑN$(�� 