BZh91AY&SY�(#� �_�Px����������`x��.��@4A@�V��w�1  ��M1F�IК h4��4 �x�)Q�L&&L&�40��`� �`�2��i��I4��0�cQ�M0L&L&T�C@4�Ѡ2h  E �	�4ɤ�7��=M�2=M�=�1�P e�v �0 Bʠ���Eg���o�
��D"�@U!��q�W�E@�T����Ro�É�3�Ͽ�����`          �����                    �@ �   L̟=�nUw�{�Ӓ���&<N)��k��g��D��Sґo3<`T�+6��p��7�UQ�|n�U�E�%���L�d�!MJ�A�
�	���w"D0�ˑ/�jP9�<��LX33	����F��S��*���|7Xv6�A��Ǽ{�����w�v�����1V]
;sx�W7�n�F�+�w�+��O4�
�j�,�������d.|�a?;�=-��B�L_Q�h,�H$i�H;�`��'2u��ɻ�Y6�$����ZT�q��/�<��(��llڤ��hyq�d�m�LdK�Q� �1y9����ȅQ�5m��b4eh���3f�B������I��[^g0Sb{��YF��<L2��Wj"�ʕ^`�xF"�ҵUSY�5/x�J�i�ED�X�cL4����;.*�*�B.\��es"�nV\�B�����".EkR�gU ��=���7�Kʹ���t������k�DR" 3{ĮUkeHI��a�C�/��Ґ$r�g�F��ds���������}������;";�0H�q�y;�].�H�Ŋ�����(D��Æb "��ں����X���VErr�0�\�������5^�Y1�s�F�` ��?VVE�S����5<�na	!RwSт#?؋Ù��ӳ3On|�/{�xH#����tA���-��Ēx��K�m6p<�-d9�N`{5��{�ݚr��Yk� �X�!������$2Y�r��7K)Nh�2�Era�ٵ���:X{��E�9��V���.l�t���d��`�qe��n6����0�cr��� �LI�R�Dx�#��w���I`����BL�1�����S3He+QfSH��C�MՔ�	����/=5Zn)�GJ��10��Uz0l�����%��{W����iR��(��Dۅ �jXs���t6�`[
E��V����=.ZbO��*�l2t�D8T$oȐ��z��B+۳��<@�W!�z=y6�i�sُc�x;�qPӤo���چys�_�^S��Y�ѩ��Ty��X&Y�[b�B�p�tV�@ ��K�g�㉒��I�Y잙{�Y5<�i��'w/{u|�-$LBKMc�ϊ�^,佇���	a� �@�̦鯽l�F�U��wu}#0����eƐ���y��3�w2���?%G$8�����[����	q#!-��4=Hx��rK�.�Nr�E����,$��ۧ�>��.@ ��l҂F����vGhF�WnY��ʨ}"t��c#n;A	�_÷[=c�6j�@��z���vͮ�`阡��م��S�|�+pK��w$�LL���63����G!���p�xs�ʐ����{#1V &����ܻd�eơ���lIqEp�!��+���\�`UU]�y{N�y�Z*�J^-j�xl [�u�Jַ1\i�R��ώ��UĬ��`ˊ�����T�ɹ��F@M�a�a�Mv�W���@�WD��)����e躵hF��/щ� ��=ٮ6�ũvb�<d�ӛ�����M7P����\�;����+��9Z��s8鈲N����L��̋x�3[ 7w�E��������8�D�/c6B�)�N�wu��B��Z/��%V��^�t�2<��ΦQ�)�y��o�u={ذ?Q�.4Z��y^�T�[�A��{O�C�͍�QD��%��^�o�TGo-�w]��|����<���2�k�N�q��q�(���uZ�� �2����O�݇��:O�HGpL�qx/�_cE#v"�!�7|�%��W;��K�0#ݎ�z}U��x�/��|��祪���4S�K��Y4�ѵ�}!�$�h�;�|�Z�6"�z��_�C����Wc#K�����Ӡ�����Yf7{7� g�Efn�1�3�fj��]Ui��t��XO�6���·L�7���1�����`./IlM�z����]�."Ces�js�onfÃM��uY7����t�=\%y����S�YQ��TV����=eP�����%�gU�@�XK	�}��=Q�E�Ѡ����8e�(7�  *3q;��FV\rYI4�=Ъ*�s�@c�Z����$D��'�Dj@������o�p��w��=",Z�=�qgj�f599p�w	�o������q :a�w��{H����)�g���d������a�=Z��Sf�]� �,�������A�N�	$�T�#���F��>%AT��t�YP�|�i2��G_����GF��Y�Mӧ%���S�;��$�QEjIr��,L�"9n�<��≑�Ɲ*�U&Evs[B
��s[C��DӰ��Wbq�5�1��,bv�h�2���I�ƜI�¹�ǑqE�DPY�H����s��2I׷E;.*��,H�����J����,:A��At�=�n'Qd�4����I�tYP\�� �r� �� �&����O�{�{��Ċ=�.<�����}�ܕ=FT<����k)5����Wk��M}�r3ES�t_��xg{���?A�ES ��b	�h9Ǔ�6��{֒O����HU��/�7c<U�R��T-�UM7O|,��,D�8wY�H���)�n�u��||v=V�؝i&���cǮa �
:v���Up�l��QeDD0(
dE�\��(;9A*dwP�r���7B�+#�`��+�����#�1���&bPOE�DA#(De?3aw��6����XG^[�[� �Fa`U>v+��0�g��T�S �z�ӕy9l�Џ-�=�<�����z�v738�>�πs�Y<N�xx[�MT*�X���ky�m��82��v�����3�S��}�	��61)ٗ8��d
��*�����V���>�V
�pA��A�z\k&��".�|�JP"�"�I�����#���;�g�y`U"�^o�e#n��
�vz�)ώ�J 9�A�y�p=叮$C��&�f��8h5p뼏�P��#y����	"��*�`���N�U6T�S�����x�m])tA;��!6�B1;g.�8��wٹ�ilN��&�s%�c׀*��:��3;]��"F%�0�ӆt�_|
����"aQ��Q3􌺡!O�gxL��kS�]�-�T�7�L(o�'�Z�'�m+h/��:J@�S-#�rE8P��(#�