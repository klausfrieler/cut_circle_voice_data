BZh91AY&SY��oh _�Px����������`	o��   ^�@�($�M4MQ�6������=z��4H5= ��  @   �0`��`ѐ��&��OE*        0`��`ѐ��&��D�Ѣ	���OMC z�z��G�[\D�nRI!IDАp���q��eM��"b jx���|f� �i#���$ ��T���Z�.u��^�a�d�9�t�7%������3fE��ݭ�]��]�T�_��!HCO䨓�L���롖�(!K�Vdzv���U�ī+��LL�QR�rF(Np �T���"ڲ^���GT2�%����S���4�Xo�����>W�?�7:� ��v��H��Qޠ��)�
0��OD\Q��Y��X{�i�$*���jԅ�O�,�I$�7�0H�G���g�ҵ3���%I��Ò��5��s�R�г,�	��EY �}�w�+V�}0�5s��U��6p �¥�Gr��N�-ǈV'wv��<	f�t�a��3 ��T��$�`~����zm
�<)�1+>��u� /{�r�=�q}C �%@�)B�A@-S�T���<�.aF��A uA$a�Ka�q�u�?,�  �)���҇au2��wL5���l{q��@�\#�(���C�wT*U�[�d �ܧ�9�K�W�qR��3�F���P�z^���X`B�"'�^���y}TH/	v���4=�Σ��`�V�T=ݔcL���ДD%��c�%�P�Ue�>���&r���$������PY~T�(P���"��E�P(����FCB��5��/&�Quk'	���C��Wd��yF)�g���z;WjN5)���	���l�Hк�J�Y�-T�Q4wL`��*��W� �TK���*�4�ɻ��2�AT
%����y�Z���F8��d�g��1�$V�Hr�`>":�[v��4���TR�A���rƜčk4��6,�\#54@�k���7�A�PSUZ�}���nH�fbmE�B{k�I�;��&�g(=Fd!wW�I%�b4#�V�κh*�O1U��.6H</}�)*����0M�Y���;�GE�*����-��.�I�[  Ի��)[�����s&o G Ո)��ʘ�+���_q��^��		=�H� ��R��Ws7�( 	VWJ���~{�"n�K(A�M�P�	����
L��*Pl��$�h�m ��(��]�1fm�14��5CSt4�q� ����4 � $�j��Q�
/d��Du@ԘA�X�v��V�y4\5�3{�f ̐&bl�s�l��馏9L���m���p���������iO2�EM�ý���)Ȣ��@�q��[�[�v��Ȑe9�9)]@w@8��*I�oI��f:_�z��w'��#��M�#�z�{,��Iw��Q��-��MDf���5�)/,`��B�U���#ƽ�`��.��� {�Ǒj���I���u��H�i���m!CB!��*�%����AЂ�VJq=�z��;b�=d���=����ژ������+A������Ԃ� �N�"g�yhLi F��Ij�E�Wvu���9-�W�Fj&#����3����s[C�(�o8[oey���Ѐc��?Mi��K�^^w��լ 9�,@�[��໒h��5� 5ȹX8�" ���,�&�&�;O�c�D�Z�f2A�Iu�i$�a@��"��6�/Z�Ap�SU�SP��Ti�L��T@l���Cס� m>2	jʲ����#vٛ��p��x�encF�k�􆦑�A�5��:�	 ad�	�K�� � �'O���5u-�c�E�6:	�8	)����F�oRkfݙ,�$V�=)��JD=�[� V�М���1fg��A�>OA}��J�H(+}���SC$ܛ�y�R�-�$nU)$�KR@L��Δm��g�����3� RF]�Eo�]��BCە��