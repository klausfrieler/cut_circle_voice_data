BZh91AY&SY�$t� %߀Px����������`^Xp7��d%!@"��(��HD��� �|ۋ�R$$��jj~�<��COD�@�� ��ER�a0�40�L���T� �ST�4dɑ�aC�M0�*R��H� �   %B!��h�4  h4d�MOAS���&��j~������i�b�E%�@iD+��*��U+O�
ԸaZ,�R����g��T��*2H�d���D��Yv�kl{!��:��^VI$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I%��F������I$�In�����Q
RJ�"P�� m�|�ĸ���&>��L:�@|!W����V�`�Vrm�S��rݒ 4�yy��؆�����-Gm9
��.�s)yu��i᫱�3�
˶�t*�~i����/<���#�a8f��cL��N�oN�U�:mU��e��f�Y��u0��42+���L�ͽ/�FޗK�N�xT^[��Fs�i<�i��F�_��fۼ�1+,u�]��ȯ�$||��� W{���>Cy�U��U�����bظ�,T�o/M�R�X��"ffg�V�6�<�;�v��j��9��vɺ6�&�,-���Xe{��ό���;���D[�**oO�ۥɎ�ej�Z�ϛ3�m�D���l�	y�Q�T����Z�ur�ѫE�`�� �o����l�R�9(f<Yʂ�<Pm$6���:�%aYJ��Fz�bqH`a��:3+	g�y�|�kZֵ�tU��uH0v�����0��+ý
�5'f`��y���	n�@0���ߕR�����z��C6nky��Jk�ڻ���:���!�zZ��n�=(j3�7#"�[���ךp��#W�vi�%t�]�Ȧ���r.AYx�[w{�|n���6*�^l3cԷ��qdLfgۅd�}ߴG`X��)����]T�yCE��Z�������A-ߔzZ������X{�r�O�#�H��}�� E&�gù����z�}����ؒJ�Z�zC#�ӈ��4��#�p��WK��a�k� �05�	 ���i 9�����z���z=�<e�qf�p_��i���|����⽯_7����b+Kmty������xOƿ��?ի9%����
CU�꽱ltњ������ѐ4�"����v5l<�1�OG��ُ�Ot�����z;x<�������}jX1ņ�����(��2}a�z�l�>�����yv�;,������Biox�I�|$�5k�p���Q@���vH�8���0O[�zt�6�0��3���>��CP��oc�m�v�H���TH`8 h����{��vj�g%;l����m���vw�(NMc��������"�C;�g��z���;e⡱bQ�U�$��F��p��ew����2�M5�|��I ���,Z���W��r%���\Ks=)�X-lBK�Q�o ��"y �c���&�F
eP�8{C�O��>I.�Ӥ�f7�W�Ҍ�tLY|�d��\�p"�%����/��S�e���}��f3��������(V�~�E��b�},Tl�n����R޺�~�Q&+��M�U��M��S� 5��hw~���+Ό���-��U]_T�V��\0;Ņݾ��*dH8^�kC�<4^������ab�弒Iv�N^(Ң4J�lC+���r$�Jd��Є�,ћ+=49���>��r��զ��t+,Ec[�ʎ�،33F����jUoJ!*����ӳ��&c29=��x7�c{"yN�=3�%���aV1X5���;�DpB���d0"����$��z�L^�jI%��Hn|�c��j�*¥�	/���������1#mt��g	1�.�	 sqz3d(���R�������} ���=���$kyw=ؘ������ <��0�o�OM�5Ѩ����w�������q�l���2#dp�Z}��+�WS���9$�Z����'���hfI���R��Y{��kX6�Q���A��M�R�7U0�'��(B&r��b�����Q�i��O�˰��׌��CU��sw�����^{Gcmв�&��[x�5��<vCsD�k�֜5�}���\�I.��\��ڥGcU�L����A��^Q>)u0A߹ZpzU�g���!]c~DuhϏQ�m�(lc��4t��Q�UCp�q�E$�c=������4Gܥ632$�؎�bA�o;��*05K�;�n�olEa~�] FB�\�\�;�޾a:{�FgU�ٻ�.TB�j䬷����Uit�Q]�42��L��/F���V���t�2n��A#΄U(�����x�.ǄC#��&�-�Rr�3'b�]����d�[�ŗ��:h��qm=��)p��?��$�A$��HJ<|����C�Ĳ���m�(!�V1maD G��Y0ل����Q�)$�5.�u�9E�$� ��\E
�
9I��rH������2��ea\� 59G9&�A;��8�m9�P3�n:S�s�)I&���!�9�9CA&���D�s��%E9)]�t�;s�@�tK1b+j9�Np�q�&r��!2�2̲"�Z�Ap�<Z�+��S��F�^��{]1�wW�q�\�|� 2$�QΔ�r}����c}s�|�O���j~�׌-N�ܠf�o4��C����P��N'���F5꧂�zmA	��ur�j� |����=�k!@\�bo�M7�3R��<��!T�FۂZ�.[Vꂘ٩��$0JY5��)�xE���1*V={�G���,	�yJtS�@���жQ��%Q�Mr�w��xꈦ\�D�T˲���!.��A¢�˶Q3�P"8۶ lGk� I�:a��͊1�w���7�{y�
�Ģ�,�����W�kf̽%�{�`�Zp������\�լL1�Ra�	�8w[;��XtmQ�����e�$j��u7��č���c�x����]�ܐ$dla!!�������!��kT��w.��yM�"�}�<:�剖<niJ=M�a�4PR��L��(>H��i�ǶfY���Ҫ�r
����P�,&�ԥ)I@���܆�����t��0�<�#-Xc1.����=��9�Sz�����G_�`$�`��s���(}��,��<�fդ�����ğ(sE;J��A�S,��a�ԞU7�

o���x���37����,�6a�&8�.Qh�s|{m�ۊƐE.n��SP������$RWԚ&���nL�Ʉ�v�:�Ր���B�@$+�HF>SNh�O���O8T�q�l���b��ۂ)�^`E2���G�kH�����C���h�~��o�]��BB��҈