BZh91AY&SY{� ߀Px����������`z��P��   �8 � 4�C'�E4�&z���6�h =@4 jx���Q��	�� � �0&�� �`�2��I�iM      `�1 �&	�!��L��R&�4 MO	�G�&�LF�G����K�A>;D��`(Z ��ʥq���'�4dU$ f��	?Y�-!S�d
�\��>hä�V��8����I$�I$�I$�I$�Ia$��I$�I%���I+���E$�K()������՟9�w��F��[��9L��aG�}�n�G��_/�1Y�c�Q5�����0�^��.��b��u)�g)��y7��5��\���5��fVEV{OP��s���Y+j(#"�v��� =����sf�D�ODV�F�M��Ys�e��\��q�wkX�r����S��W?��~�؈ڮ���#�F6	�n��,"�m=cBzee�ٰn��;��6��m��9VP�@��&��ܘ҄�-��Ʊ�tr d[S(���e`���B�w��B�ff�T=�f�<�k�Ÿ��;h^72F���afa��(B0�$:�IN��f�w��f����T�Ph[�5F�J�E����� ��Ǒ�z޷��r��0���k� H�5c]�@�w����(3FWA�	�d�@!�}��Uᇥv�r?yB�E��BL�F�;�=x�C׎`D���''��dM�zg���T���Eg)%j�Ԫ�l9��Nr�Wxp�����(���dyU6"��y=A� ���ǲn��&�9Dof�È� ��������t0��>�g��m�]Q|mV��K0��}���<���/\��x-v�"8*z�ח%�����d*�.,���xZε��h���]�j�"^}��o{�9te�; ��;p��U`�mt�f>I�x�1�o��|�8n�dѢ�" �a�2YK�h
�������hKA\i���t��2G�����e�c��c��'*O8�<��y�Ch�H�`2 �OO�����h��	�3�4���an����kU�U<�_�'�X{u�{�h�Ъ	u]*�P�@^/�	�����8��g�fiGC���^��L�$�/6���@��݂�O����C����� �;�s�;/TS�R�mc�pU��X�c�q�����0�3�.aO0���#N�	f�kww�=W}����R&�VZ���OD
B�`��G���q�'��0EW�^������Z{�;�.WhS2 �n�Q禘֞ʥ�i�W<B����0O�CO����@������&2nk ��ܴ2{yæ��s�����]�+���T����3FT�����E��� �W$�>��XGE��Y���E����ǧ-GԜ��VttE7y5�n=B�ׂ�1�* {������X,D	*;�I�+��s�E����K�q<}��S�X]�=���r��5;��gם����og}�v�:�&���͓!M��^Lq�Fިܜ���͟����ק���SqEeҔ52R����l��ˈFJ�=��ܡ`�V�Ǒ��*c��ѣ�=x�uͰ� .�YS���pc7_ӽ�0��؟g����ogVO�:V�{��ș{a�'m!I���Fr��c���J"����w��ĉyz<�:�hߒy���͆���&{�f]p��:�n� Dxv'��]�3���ff��,m�B��o|�l>�5V�\�\���{����[�z�X��c�j�\!����{q�\�D�>G{�Ý�t��:C��MUi���(܇d(kS>��^/c�$�.�\�.;P�M�u'��v�,�=[�����������QW���� R��Y�9���N�d��f4��˿����Y�e��L!�Z�G�[��[akR�e�8����i���D͵(�"���*����V#-�++ �-��h
0�d#iR�*U����+�F�UJ(�-�*�X�[�`1e��M���e��QV&�J�1lB�F(ګ�ڕ�kI��5N3���l�M�1�B$0fbB-N�����<��3<W���q���|�{�_=�����97>��G��zJe"*�.?���t�3c��@>N;r�xZ� �T!�(� F�$a����Ӈ���d�}�E����������=��]�3���Q%Zf���{�f�2^$���c��K����H�)]�u���ٝ�dp�ҩ5T�u��t�+�"L�bA" �"�)��`���,� 1dH�U���Q��9i4d�4�Z��v&������MC;�9��0n� �H�0��O��W�Vf彥1���ыXfo$53 񰧧0���(�2�n���N,�����U���Q2�p�#�V҆�f�g��0�p�'q����ڈ3D �X{c륏V"}Zn�Ӻ\:�! �f�	�� ��}	u�v蔃L��ì1";J%��$8@���Hc��^Q���b�o*��Ш("��̔��
񓢴6l��Zsc*g0�j1�	��k �-5�Hӕ3�z���#�D' �;�n=Ň�$C��&�&i�6c2�贏Hh�9�5���9�B�]z�X!x���@3�H�g�������/u����G"WE���6�phu��#�k�z����&���CZ��U^$��,��Y�0<�2N�q"�o�ve-� �RvH�Po��L<��H��2gHL��fD�L�킀c��P�5��JD'��R�<.~pl �)�L^|�w�.�p�  ��4