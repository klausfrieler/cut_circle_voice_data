BZh91AY&SY�v*� �߀Px����������`�|�@:h >�   ] �^�]D���	 �&�	�L#M=A�@ �� 	J"@4�@dh�  i��& �4d40	�10�I)�OJ& hhh�F�M 6�4�=��0@�4    6��"�M& ���f��d i���j�]�V\��&�)�@ ���$`ej,mIN!&i|A��9Ā$�y� �LI�����{Z�|8�L�)K3�7wwwww4���������������ݽ�u�����;��3.lV����ݍ���ݝs?�kd�?.%�C�ܯq��7{���le*�0�\z�-���w��yF�m'W(:��ȋ�/�Oa�Q��pAE��g`�	p��`�[��EMfL�	�����i�a��`\���]�;
��T©4T�=��jՈĦ,۴�O���ϺI�O�?��gϴ-B~߂|	kV�}�/�e���ѯ��}��� ^�2K�h���C��=����Rg,��9��JWuP��Vl=��^|╈���1P��*����cAm8h�W�>�R^J_e���!I�}�|�u�u	@�on�=XNe�L,Nշ�2q˫��s���]�����BL`�Ò{��A���a<+���g?���h��a�s'��^��|(�|�������7no��o^a��l�+�X��s�+���׊��ݦ�è
u���I�)�ſ(���]�8[z���Pq�#F���k��=k�]vq�e(h�w��e��3QD^�F�Ik�tZ��wވ"PR��L�?l0�ArМ��w>,t ߪ���`��Q<�]��E&`P��Y/t� Qm�sY��uo���~��]3�#1���Aj,�hA@z�}'��xJ��ە����U����v��O_��4�25˸��ϣ�x�!� Ґ�M��g$�y��Ň49�Ŝ鳗, A���m� �b:2t
�a�|�n,=�OYʌ��;"�4l�M�@-�4�O�i���|�x;m�O��=�=��ˌZ�q�3����Wa���Q��j��+��% �ub����"<��F�C�i+1�H�ؕ;^<�E�Ĩ_�F2���<��a�23��#�m8WezGQj�z�����C�ѩ���K�UP)E����wNo��;c�Ȁx�����/0���U�S(+��@�����Sx�W���8��Sy��Ybd��p>�%Ɂ�9Y�I��E
zy��� ��qGe{^j*�7�C��5���!�9�8{"!I���A�ĭk�v�S�^���WY�W��*W�?=w|=�d�p�Oˣ
=@���������X�5Bn(��.���k�b}m&C��[[��p���6�q�ջʉPmM�zȨ���	$���k�I8�ӓ�;`��l�
ێ�n���������@A�x8��4�û�����&U�O�z;��N{�;o�7���TGI�
��]a���b�D��}���}�^7y\���9h���+f��[�� ��l�G��v�vs{��9����#�;�.��ϱs{�η����%�GT\��!���ȱ���������2��r�}7�|��/�21�:h��B����/MK>@�<vQ�����uX�MO���}M̥]woh��Q��:�9UQ���h�¬j36΃�z]�KmuI��lC�V���n�W���q��Ǯ{��0<st7Uz<ؤ� X��ϑ�>|π|����ۦ��}�#�{��3^���(�+좨$E�#���������Qv�ӭeB�Ѳ�)1�T�Xi��M8ɉ*F+�r�d�թ"�6�[�!�$��V#iDc+*���,QKJ�)[aXE���lr�+V[j(ѵ+i�q�RЪ6�V�-ˆPC����3�c�̥���-Q��5�V�Z**UeU��liB��UX�f��EmR�h�jl����HBl�VB�:�䮞������)���;������J&OE2O�Q���O�)�%2>�챬f9*�;��.��~�ە��0�\W�lX�A���B�3]��:S�G���4l_��ǵ��[�V^m�8���A_`���9��I��~ϟ����J@2�*��7\���n�u����5��|;u;}�
(EA���"�P-�Ƞ +"�X, ��� u�9$�r�v��]��%N܎�,���L��"�bƐ'R���L�W�Qz�>;t*�Af��ȋ�b�z��2���-l��Mqw����ܹԇј��rMn(FJf#K���PgQ6;&;����j�m�O-Z���8�	&:��ݙ>���9�pe���`�j1`$�u�	um])4f�u�dJA֙s�nQw�L��$9@�֌�C��X+��3@@@M��d ��amI �g������zu�*kP��c���xBGI��ww�z��I��$��f	+� ��<S:ʎ����7��M�M<u��M#���kż�6��SP�0��ZB\Jq.Ere�Q�6�Q�S^����&m�@,�9�\a��Zϧ=�ꢊ�5QE���z�gЄ��̉ĸֳ�w�Č�a�ћ*i/�9Y�D£�D˦1�	����g L��jD_J�8 Aj�ί����.�uF���OF�&m���)����rE8P��v*�