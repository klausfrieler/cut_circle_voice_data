BZh91AY&SY&@' �߀Px����������`�,E= �P �  `Ȱ�M4�	$L��ji�4!�=CM hh 4OMQQ*�M2Hɐ �ѡ�& �4d40	�10�I!4R �=@  � s F	�0M`�L"Q4&�FM4����'꟪=OD���F�~Tz&W !=��"TF�T1TC��Z��j��Y$EB�P#H��˕��82Rd!Nr��>��^���庾gW�m�z�m��m��m���m�m���nm����m��m�ۆ�m�l��m�����[m~߀2H����P����&Yﳿ ������(T��̳��9F�M�� Fќ�w��lQZ'brIUb��]��黜ɹ�a_��׹��p�s�
�n6�@���Y��!uN���H�nfQ�r	�LU®b�U����kNo5P���Db�by��d�F�LNW�A~�36:�� �,0qV�f����1f/D�-P�#��ȵrR�n�:��Z�ܙ�dꛒh���UdU�Yy�b"mκ��9�L�S��d���)��"N��rFQ� T��#*:��J��]G�}Cӆ�ua�2c!HlP��ܤλ�H�r�Q�v���B�F�u�9)9Hf$\\�Ӽ��r�%6��o���H ���ςv���6��?O��~�ʹ��G>��Q� XjE�E)�����6n*���kM�F52�(2H۰Z>�_^~����2��J�=��S����ˬ�\��FuZ����GsiK�Eî^wGL���7�L��i�:v�T�ྋ����xsr�n1�Ǫ��;���7[~�yk%a��ٟg��o�{��ʿ�2��9�xH,��k��	��w:�V�O/8��~�}'.ɳH�n��i�ɢ��Al�P��J� =q@���_��_{z'����,��$�	� F؅5#��Bz�ޱB*C����й�)�����+_;����p�jb��q9���ZyrA�j�L�̛)ap&cgG;0ǣ�Ow�D� � A�"<}��]	܋�I�A�=p^�<�kR�BuE;Q`@ޠ�0�Da1h��Fݐ㐣���g���	��8���A��O�x<�	Ip�ܡ2r56ʧ&��r�ޅޮ�"��iJ&�����}��[�F�t��OS\w�zs2�^�Og��q�s�S�qө�`����x�=��Ez]�
�r}Z�7U���|PNo����4�6f/�Ђ��)�3��p��\�����,�pm^�B[�N&{�?{��
��'VM�H�¹�#L�`��G��b;�x��ϟ;~�:�Ȱ�=���tc�6@������:�v�m��u4Ñ�3��Y:&��ی�����BQ�DT�,9ȵ���0�cL�c����:2rI�mF�!@TP�xN-�p�oϽ�c�̧�R��|p(�!�)T.0x��������쇶U��:I�Vy�����l����Xg�1g��=ƈ��ՎVn�{�Vi��{7ޔؚ.��q#ٙ�R4k+��W����{޴��c��2�sF'��1��څ��ɖ�"�(�=>����H8��R�"��\���S�LgfO`�tA�$��Ү�` ��s9�z�n6t���yr�;|`��Fxdԥ�7{���苢Կqo�����DcĔf@���wp�!��7��F�M�@�Iґ
cϝ��=˛^�]=�M��Զ����3�<�n���z7cw�K�:�j;}#EԀ�2���7�H���F�!�3�{7�s�-U�w�~�{�+;��ٹ]ݚ�j�������V��� �����"��������ӹ7�2���ng����艙�s2qu�]]O�v�q�	MzD��{u ��F��E>�_�x��7Pc~�^�V�#�!t���}ЊQ�v��K��MW���4V�݉�7�[�a�)v��
W� Y�I׊jD���V}�^��y�
�ݧud&�x��t!�[��4�BBI�	$�
|oiձ��� �o�mti�w����|�jұ��0�A�f*1AKJ��XTYBQ��)1��U���T�  ��6�,ь`���
���E#�ݚŚm*5�PRԶڧ6c�J�Pntѥb�K0b��2Lfe.�kA�0���F�b��UQb�5*�ER�[q���e1�J�QEjUUk��ғ�q�x��0��<K�憏I�* �f�T���꧛�%r��8]�@�Y��/�ӭ�WiO24��&�����S�UU�ٕ��a|����m-B@v+��xs�Z����?aފHFՐ�p������l�ҔO��gP[�6myN����A@�JtC�T�%,�*l�k=qj����c�����w�\`���эRUT	�N��4�S>0r��yݿ^����u�AI��(DAT�`�
FD`"$E�
(1��1X�p2@�Xl�a�<,G]���f��*��k�i�wu4
�T*��!��|����ZXj1�-�󮐞m��Ƞ`��0����?���0�HfN��726�j�.*x3��[涑E�LF�᎒&)��c[�7Z��e4s�H$�fI im�Λ���3�u�X�oB�&PB�P(�ܱ3c� �)@�R� ���Wɘr��"�k�s�p�2,��w�H8!��s�2�`��0��	W�G��/[�0��Ɛ��ρj���(�bl�`��К�@��ar���Y-{�����H�3�W-�97=͢���������>M��xB��f�]�"��'`(��P5X���0�sdd����Η�4D�̓�����5=ژ֞�ڭ��*cI�ڧNY�@J4�=�i�\9cs8�P<6d�����@\E�p����"-�k32	���OT�q�i�mNN�h�Ҋk��tyZ�'��[q����C}(�,�x��rE8P�&@'