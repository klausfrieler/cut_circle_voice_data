BZh91AY&SYa�) _�Px����������`	~�p�k��  �*�TP�SL��'��b�LL�h 2OA���?JdѠ�hm 2h � s F	�0M`�L4�yb4�d2d����#@h ڪ=      �  $H"i�!�O�O5A�=F�4z��G�?iI�s@�$!؄'��������(�m��P��O�K�4��I��Y!,�I��������l�-�i9�s���333330fcfffe����[����w�����q��qG�?1�=�^y�"u�x�_I��CPr�4dUL�˚M,[�v�np $�ͻ���F�dT޶�Z��no2&V��̸��\��q�_��<;�LLV�{Jh�2G�t=}\�_`��^VT�^e>U�w!�
�Xb��)����[@�R|"6��8�,\�FE�������u�6�_	A�N����rf�)�=7&�$\9u0����F� 1���K5��S��*Uw�B� ,�R�<'`�,&��D=��7#��n����U1&�XÚ����s�5)+�cQ\b��6�݆����Uq��#�iu��h�Á�3/d��1s.�b8์k�}#�x�a�$O������Öb��|̚�Z�]���f&�d�uok��C�8}��vpv�}fy��(�z �nY���.q�i�a�7���B�!��Z��ء㫺~�#���yv����N[��*���uv�k:fpC�9��v��+��N6qTB�]m�N�Ys��E�ewǗ�ɥ-Ă�:\��E2y���qa-L��[����Ͷ��SoƊ���c�1]8��v���-��N&��ª&f���eֽ5rzҊ��s"��������iNMϚ�e!����3f1�L�E 6��p��;r�҈9"\jz��\&{�}l��Py�� T4�m�5ơP�����:j�U���쮲�l�9��f�B=��Χ�˾��x���I�ȼ����D��JYK�1�ti����4�ا�h�t�-�uB��5�f�tX,������0Ya�<L��.�k=:�@z�N�_��Kjr^1R��!�ⰵ�+-���Rt��3L�����wz����Am�'e=��h�ֱ;����<\�:8�9�܌�WN�M)ѐ�e[q�M-�lm�1���/�{{{6�( 	ZU�)&�휉�:�f1,��.�H	YB�Q�/��`��$�����29�� BaZTX�fe��V
� #l�dV��F&b�o-ݑ#����"�,B#!
� ��V�q��f��h�����n`�	��*Ye[7U��)(֞<k̭>7[^��˷�ӎVjN35��������)ąB��ٓ�1��O��^�b����������(���I��3oؽYy�;�ЈG���BD���/��jK��-���s6�4E�F����iI|1�D�5�e�|�#��&�DJVʵۆ�U�ϥʓ�9�Wep�� h�C66��"B��+��F
E �A	�x�YfJq>�=Y`���a#b �BCjI�3& gs�ϊc"\c��M�B����X@lS�@���.DƐiPĖ����j쳫F���-�ZǣLG��3�gN8W�-�הb�����n� f4� �{_���bK�U��pf=]�P@t��D�w��}��\@j�U�oD+�"�Y�M 
MFv��ׁD�aPf2A�IvT�I���DC@6^�Zj���MZ�lMC'4ea�I2�qa 9��_U��Dr��wH�۝gI��=N��ǋ��˨F��D���rl�Pii�Ƽ:��pB@�%Ęd���� �� d���#��Z0��Ί�:	����ǁ�(�f�&��g�_"45=�('8���M3_L8��U,Y�� Ӿ�	I�Q��#�_��o2 �ۇ�
L# y^?%E�3IiH���B�J6�q������{��3� ċ�q?��H�
7�� 