BZh91AY&SYym�� Y߀Px����������`�}�� hp�*���!�2��O@���Q��@4Ѧ�������@  z�  �`�1 �&	�!��L����%Oɩ bh    �A�Rb      �  ��Ҟ�i0)�j����6H�~��rh �b�@������'�m&�HP��/�KƉ0H�Wd�T�(��hbѡ��ǫ^�I�R���s�c���,g�&�e��x�Vy�������λr���y�1E�zX;����� E��)#^L�b�^q�2�#�#��;}EH���M�����47'ue;fWk��{��5������0٠X�^�T�2�BV��	Q��j��"u�Y�8�˼h�b���j:�1��Z����^��DU��iUb(^�P�6MM$�8b8���;�ԗ���:^�q�Z�-��� N����TQ�IME\�[�lJ �ʢC���8�S�A�ۈpD�U�"j\D��Tl��v<G�{Y�r�%�i⢦3���ҨbGd�zM%S5 tNg"K����ba�ګ�u�|^42j��)J��	
#e�l�㮺<^A���o��ge':�����&ﮜ�Y�h-��\)}Yd��aDI��t�\�Go�cm�P�
��tk1ӽ�F7WI�x���2y�x��6eg�DB>찬Km�̌�E���KZ�E�v�8�Y��8�y**��|+;4�컉���B mQܑ�c�E�(\�hxli�e՘�|�PjW�_�A�w�F�*%VD�صa��T+޴��/6U��.`!a $D �/�|��e�gOyQ7�Mk(��4�����m H����%H�A CM��H���!7��b���,.��B�:B�&ډd����f*�\u�+�cB��E��,�z���������u�
��u�>��O�1�By�j-T&�����J�@�o*��vc|F.��*mEiج�������<h�mH	����&a��,5�2�U���C��;kHT2N˂�k�۰It\�X��m����\��F��iJ�g��%�[�O��=��F
 ���V���eߵr]�9�!R�e��t��,$6
.4"��
J�ւs�2�E: ���L�^<	2( >"I�@Ӟ&Ҭ/�1��1M�ԕ���e��	����	��ژd�vD���lF�u,X�T��Q�rIj)E�HFf�AIzy���!���v%��<ݷ��F�w>��ܟ��ݎ8Y�_r��@��<kzL�Gts���Ja�3�TbB��h�F�kȪer�39F��WbPP*;I��Лz�rY������MC)Dj�Ӭ��q ���wH{�#h�|��;:tZ$�T�p:<�:�,ᕋP��˞��anl��#h�xׇa��HrIv&4�<� 6�ڞ���>y-��;~�f�Q3����%Q�i�^�,`����֫��	�)��=�L��B��brj:�.�E�C�LuSa�k+7��H��H��6,��H�G��,"��T�Ւ�@k�Ȑ����Z��Y�����侬g�s�lH�}�]��BA�#�