BZh91AY&SYzW�� 3_�Px����������`?,t-�PҀ   z �\\Y"��	"�	)���l)��SC�0�S�JQ�L� !�� 	��aOBdI6�FM4�#@h b!��IA4�Pb0A�&F����1C��b�LFCC �#�ɨ'�M&��bf��<Dhdz���<Ԟ���@����U G0��!���Z�n�_8^,� �e@#H0��dIp�#���  ����N�FÏ.�o�Ǖz*�I$�I$�I$�I$�I$�I$�I$�I$� �N�_�v�wwunYxu�������O�����7�.4��XD�Bj�)Ra���*2�3��ة��t#��>A5WUnl\�`����xpL��>�����W�"C�W�lϫ���@ )��;lY�]afC�O/Y4���at��^0�j�j��1R����jf�����2�2���ENA����Hj� ܸ_�"���.����1�pM"�w4o�.ʌX���q�d!��h�r��Me����?��wi
�e8��eJ��T�cƥbѣ�j�N�"=ԧp�h������8�#R;�6�6|�&���;�Дf����"�!8Q��TUD�lhhA�4�9�x������CKd=yN����V���@XP��uJ��7��J�:1.�����r�]숚���>���f����Yx`&����>i�%�h����PjO�7�0�P�vuz�ϴa���5�f%�6�SH�ц�MɰCE��;�&�+�fbU���$d=xK"E����y�����7��v3�5~Wo_x��|\�g��0A�3����|�A��F��G���玗0q�φ��C��( ��>��]Ϝ�[^��jZ�s�\ �ב	�-iL��1{N�=����#��+I�n�.{�.�M[j;��41ƻ��t�ӷ��ZK��m:��4����}�&���ԡU1�^�|�]u��|�̿��B�qQM�����T�I��N"]�3~2�p��k ��%�Y�,��Ar����7��Q��ޣ��Za@�9�C�v~��8@D�r�+�My1A�	�J�5�y����Q�>��6����g�o�v�l��`�z)�f�`��ք��>�%��!�MUy����w#�i���箌̃k'���<�dV@)�E��#�>G�`�:�ݢlR,'<K_qz�� s���E\�Ur�="3�y\=	,��̌�����j�
��!"=��q
�7swN�]��pY�Ɠ�W������E�]����ط��^�rB(n�����{R�u	��̷��H��Z&�y���;�6D�
"��b>~��oG0&��bc���$<��[�UTs�8�[�7���:B9�\���[���+f�[=T����Y����$����� ���I�p/�D��*z��,�q�Yf�K��˗1����{9L;#碻�e�1)���]xR0�;���5�Y����͉�4ĵ���]�P{Ȋ�@��]
w�}��<1�`	��m�C��mڨZ�p �ve�旫��=���%6����q�lĹ�uWYs�y&�}��a���V]����>���PE��2e�+��-e��΀̫�D�w�0|� r�nc:���GM�Ҡ���Y�ܱ���K���vO��É�Gu�o$�s�<?u�]Y���?;A�+3�s���"�♘"H���r}��"L�l3�-[�v�D`�&��5|]�"�1�6�Ɂ����X��2���^+���gy�Ap�&���Out��W� �0�6T��4!�3�]���ę���.��PM�KnP���MVQi�C�f� �&Y�����p�2��^�=�숬�ͩ�2�{��Q�n(}�K�<�!�:��ܗi���kA�@!֌6�8'�7�k�`�h{"���+9�ts�p����6嶟��uTE��X @(P��{|�t6m.�p�j���i�e�Z\�����aSD+�cX�մ�ţi�����kJ�h�¢0-�QB��EJ�j���RB�X��k$��`�ʢ�����-���R��8�cZ�XֱJ"#lTV[F�̥JԥKZ�V���TTNM��eJ�6֣mj-`֨c1��X�m?�T��NO��Hp͞�FUa�̶�I�I�*�wŲ�����Su�t��-^��~;RoX�A
���,S��}ڢrj�O��T.�:~
]k����@{�v��y\� ��?Q�@�G2�P:À����տ�p�f��x���
�+M|��q�:�+��T)���!d�ӆ�$S��W� ��u���������<�:)�$�o�R�nhJ.���۟s���(�K �H����`�aB�ER*H��&��:�5@"I�(0ѽ���^;��b�^�}$J� � 5dd�����L�8�0�g���>��ӽ�495 ݁~����0� �8u\ܑ�\�������]\	#9�F����H֠n z*6�z�o�Κs��8("&�<�3ټW�V|������u��P+�*�z�ŉ���J����ho*\K�pxJ��i���d]��0b�$2.��A�8Ӂtw��"/},�f[8aC��!k&�e�f&
�KC_6
M^�Ҩ��,�>̖@�A����T�(w���\}�M �=�LI�(�ICY�s�z�� g�^vy�S�P!e@4��<��=;�:�8t���i��߼p�AE�5��}�nPe�f��)c�R�MB����T�%l�@�ڱkŜ�0�oʸG2�P��	
ݒ��_��`?�t�:���	�P�����^ 3���Gu�"~&��B���(r��R���o�]��BA�^��