BZh91AY&SYW"�~ 	i߀Px����������`�p/mt    ���[H���"�jz��=�	�z�����7��jz��Jhh � 4  	�hLBi��   �MyJ���14bi�b0�4d�aT �ѩ�@�  M �@4(A4��& ��@��@ ��
�s�0i���)U�A��2��뺯d.�$��`T� }�?k�e@qH�ңBd �5��d��o�Ï.���Zֵ�j�I$�I$�I$�I$�I$�I$�I$�I$�I/����4�3�����Bcؼ�{z/^æ��Y�r��(�&,[���.�"�@̙.`b®�1vǧx�D�p�<�9۰�eL����tܒ�*��kv��WLr�����	Xe#�*�E��ӳB��6����%[r!�	�;��!Bx��{��,� ��ã+	�
��*) �H 8�,	��3v]�(ðO4���n���O�rFL�PvҲ��{�a��l��qr'+*b`]DLx�DUE�s]:���2e�e%1����+VV_���5�T�N}X�;m��g�v���k8{�ߒ@�8
��oq5��4D�F���H{�����Kʆ�[Ɂ��w�fs8HN$��U(uW��;!��K�:�'M��P��Gɻ�[Ը�u<���,NMڿ��~�th�d7a�k~q��Sqr[�8Z��S�N$8 y1�>�h�4	�k�~T�l��(��F�<���a5�)�����O{c�����-?+�^���78�>���ԩ�/�La�����c�U��V��u\w5ĺ~6���䰪�0z�T>c��-j%�-�+�|#^�a�8#]Z�q�
�C��y}�=��܍��f"�5������Y%��Gd��,�V�	������M_;�g]���cCWl�
6.�I��p�s��V�L�l��(�c8E���ǈu��.���ꮥ�Mw�o2��	��`�H�z���a�t&&f����[y��@諉zw"���D����6Af�q?H����n�/[mȆx_w���*���FW^:1��θ��I����2"2�Yx�׼����=E�g9 -X�x�l���;Mw�d_m����f�f.I2��*v`ja$Ln�,�.���V>=�v"�GA �`�xm�Q��ye��:��@�0����]�M�}���]��.ȥ}���KV>Mx,�h���.�;w�F^ĵN�osm�g7���̿d�Y�X(��'q�8�-O@�n%�&9�<-�ul;�B�Y�j���O����~�d>���T�-��5��L�1n��0=��--m��КN��o��@� ������m�����Y��aFy� �m��'�F�f8��{��:���N�ڑP�ul4�Hn.Sc��u>#i�[JA<V4��l�����#���9/��3D8��e�vb_-�ރOx�SE�\y�*�'�dydYu�y���������ùz͛W�V���̄��J��(%FxR0��HA	�*$��P�F��)j�V�{.5P�IAHaw!V4 !��n�b��OIM��X�a	���,����aw��21!�J	����+ PP��HUR"DH�
�}]�����P�u�d�7�h���~����l�V��|��h���L-�e�E#�X}.����Ӳ�&.Oe�O�C���W+UhYlK$�dt�M=�|��^��Z�]�.Zz@�0aR��/� D6³^��s����E1�7BhGB���k�oIt�L����l�!4acH�{���n�$J}/.�#T�M c3�E-�5\�]�&��֣k���ݨ^"����Y� 1'�&;.�FFP����[,�V��E�S� U����R*��9�������v�кn��E�C T�B~Y	���ҘВ!�@<H�]��>*��ԇ��K�w�q&�6TF��>�fj&�'��ߴ9_��|)�	#SI$1����\G�Uk��˸��A@�4A@k�
�</�bfǗ ���mT��9C8*W���Aֈ�u�lFr�L��]�����WU您X.
��ԥ)d]�мql��4�����V�LRZ�|X)6�I�&�t����@
��=�ʞe��k�F�FQ�ہ�swx�f)�P�#��j8B���%x�E��M�T�M7����;c�9=;	|���Á �"��;Mц�oQk=�ޯ�QKN���b�H=շ�$�N�)ļܰ �����"1���h�Ē0'@�LV��ښFF6E���
����54��rsQR�6m��9����N��U�3h�@$����w$S�	r-��