BZh91AY&SY�*E V߀Px����������`	,u   ����hZi$$P�ڙSɚ&ji�(�OPd ���S�IT�446�@ i��@ S����       $�R5M        s F	�0M`�L"�L� E?Q��T��4�$z�0#�&\�������p�<�Z+?�mf�AXX��D� C(��) �q����LI���F��f���T��ײ�믌�9����`�������������������������,0���%���x�%���H44B�ob"&���\i�,�e��"��w���s��qR��B��z����"B��swI<��ૌ���j��������C������O1�(1��("#�S�'"H@1'1J�|��Yc!�&^�k�wF�kQ�����8 ��Pm��)�?^̵�x�r�}��^)���c�5�� ��۠�g0�)^4a2���Έ@A^��$Ƚi�,��	h��&��.jƉr��}rƵ���-�>��.�������ʿ���3TD�����kO�F�f;U
�!3�C�����(w�z���C x���jM��*J�x묹��;�x�C�J\����0�䛗����f�B��"i�s�"끧��*�=�x�D���x�|o�nճ�.�m/cS#35!��k�^�"|�e��xOx�ذ���u�����
�ǐ��n�0��0��n��i��Ϭ�6�9�&��t@������e�p1택���'�� ǭn��c�L2a�6n
Bwq{A�׬��p�	��C`�"� ܭ�i�N��Wi��]�y��,8 Ԯ������i�Y@b�;�C�W�9c��-��v�{w�����(��	y xM�`�����ZA+
��6\T��cu�H.2��I���)�1�]B�C����q��U���m�xA�����דظ/"�����5Cht���ǐ��&*�$J0;:��XE�F]� =BwtP=�,ۘ�t�-A���N	��`�I�LL����OrH
W���i��eU�1E�[2��U-<�հܒ��ɧc�`w�m��x�K����gGmY�rhN:�YS��Ք�og�)m�S<gVH�̤�	c"�(�ز4w��}A(�9����Y��λ.���*w-���SG;����lm�cm��k�͝oe��88 jih������1A��q�8��R)��V[Hh�4
�~�˥E����I�h��vܖ��*�+-���r�+����#[F�es,�
̍��@��)��JC��I�Mv��f�՛^�7S���M���[S�-~�ypS��U�ݎ�
G���5��.�i$�I-
ƨ��c�8�N�G]���a�]����A��z]7��3����zG��b"�����M��{�\��,lI'a��I�!�����zK�cF&w\�d�
l�Ч)�B�������z�q){��)�p�SJy��Y*z\h������X�T��ġ�@dU�0m$5�����E)Ёb;7���f�Nm?��JxW�ad���$��M��Q�r�v5��B�^����plq$h�,��+�`��+1&1 !�@6�Y5�U�K��Ӕ�������Fw�v����'�����C
��~��!i�������r��	�+���umYB���H#��e�&��n�/p�e�J�n�w*��Hs�@�j�<\#�� M�C�d��8�@�6�nam`D*��L�nѵ�w�e(�؆+8/,�H.n貑˭6�sxJ)����"F����*:��Z�f�1�=�,����N��=[Γ�$(1W{.���D�D@�S���[��&.��?����*0s�	�T��3La����v{�VUU3EaT�ă�\�kB�'�8�U�ָ)�7��%���������Gʢg���! P>�p&~3[xb ~5+�Ű�i��((n�I���e(���ٯ�9Fm�kH�~1O�.�p�!xT"�