BZh91AY&SY�p� 	;߀Px����������`
�,
V� Ҁ��UA ��$���M14�42zL 4�����J��0� � ��M �4��4ڨ        JzIQ���MF��&���0&� �`�2��D���L�����z�H�h�@h(�L�
��y��("�H�����_�/IF�)@��?��Y@�I��� ��c.-�-v�{8#�<>/iJR��,����I$�I%�����$�I$�I$�I$�I$�K�tD1�7�\Q����xQ�ಯE����Ҫ��%�b�L�a���� =�ÓFp�D�=�8��ⱺ�����pf�Ɂ"5D��wN5ceF\�rA�/3jmb�yuMV�fp>u2���J������ A]v%�q,o#p�K���C��`��%�#́�
�L3I;��Y��z�r�AA���m�v�W䋝^��P��$ ���$eG?u��)H4!\!#��|�K.�ÿ��l��]�cYw�]�9���a�V´�#��H@������Ɖr��F��}p�V�+�BD��9��N�`����<6�6�;��DSr���E�Y�T��2����[3+G/��Ph�#�c&g%��&�e��\9<N�c�ЉeD��"�|�RE� J}� t�Y� FHz�S?��s��oDi2�4k�u��9<`H����T��n���ȋv��<�GSp?1���t�����#�q�G x�9�5��]�����ӌ�V�4Qظ�H��]ǧ�ar���uq�H�$�����v������/N��,�R�<��#���rv��^��_	S�6��8�i�a�*���v7��E����@h�w�(_<AbF�{8�ıOE�˽��ʃ�E��̜(�L�چO!��������d�0�EEc�8��gHq��8����Q灪m*��T�%�d�nV���>�DP�cK�ʨw���SY��ó�f���k<�u寂K��k�k�31sv"ZC_�"na
ʐ�k$�M-5�ՈMK�n=!�Q�_n/�#�d�#�_jZ��:�������u�-�M�e��L;L;h�Zك���]|T���$��L�a�0{m�E1lk'�3��&�GIY�Pȥa	#� .v��yvAecZӴ���<dp؀���Mn;LUͩ`&_(R�B]=YuڕL�dVի�z��*�:�Ә�{���LN]A�b$>W�(�r�]���|k�%��5��{�2�`���_��6�N��{`�a��[e�v��a5�s'�F�MvC�Hl����٥������R�m%���/�AC��g�2�<"���3,�z^v�(&�휞f����@�����:�e�/��]��9o[Y��� �ʧ��1�Ŝ��m��n�gr����'[��{#2��%	�dF���f�1��1�5�j��U����_���*"�碨5EQt�W����i5}�P��C8u��rb��B��"P�����ҙx��K��e�eܤ��q0J�!yr�UW �re[rF0b2$���E�l��QIBH܈\�H�J��#���4���@DdE�$T��F1#KJ1�nL8���P�vfA�c��1�TL膿��"�Hh�tv�K���)d�7�P>V����g���O+�'�4zPM�3��Lj�2Uy(�y_`�9'�G̛irBGZ��.׫'��`�ǭE3UO��Y
`k:[μ�v�9Sb�#�v\� �틽�U��$�B)���,�J]5���=�j��s��h����=�`Np��SR������Y����X0xa�7���I@H��,���t!F4�¶���<a�[=/ÁS2�)�dd��"�J���ܻXn2�/���О];�k�@ųP�E<1/��0�-���QJq�AW��:/����؝���^��T��4j"hO6=tf�Hp��VÂ�x��BE�fBHa�u7�tۭ��JXnbݾE��X@|�)�s����.�C�R��S0�")\���vQE/f�#;:�e�_<j(;^J�`�P�Tʥ)H��	�ǂM�q��cHZɫ2��S#��F��T��I�E'��YN�m��T�W����L�g�[Dop��ͦ�&���̑�P�G���s�SFj����ܞa�M�=�.����:��v&�~r��=A�5Mov�6'�ѧE����1�I=�]+�A	�r'��5��-�����,`I5��4*�����i�S�β�PT�r�mO���9�����j)���%�D����O��8R��)�n���rE8P��p�